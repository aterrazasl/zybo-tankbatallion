library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity M2716_rom is
    port(
        clk  : in  std_logic;
        oe_n   : in  std_logic;
        ce_n   : in  std_logic;
        addr : in  std_logic_vector(12 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end M2716_rom;

architecture behavioral of M2716_rom is
    type rom_type is array (8191 downto 0) of std_logic_vector(7 downto 0);
    signal ROM : rom_type := (
        x"7C",
        x"6C",
        x"7D",
        x"43",
        x"79",
        x"DB",
        x"0A",
        x"1E",
        x"49",
        x"09",
        x"86",
        x"41",
        x"43",
        x"45",
        x"44",
        x"3A",
        x"20",
        x"41",
        x"09",
        x"52",
        x"53",
        x"4A",
        x"09",
        x"32",
        x"30",
        x"31",
        x"50",
        x"54",
        x"53",
        x"0D",
        x"31",
        x"44",
        x"41",
        x"30",
        x"32",
        x"42",
        x"53",
        x"3A",
        x"20",
        x"41",
        x"09",
        x"52",
        x"53",
        x"4A",
        x"09",
        x"0D",
        x"35",
        x"30",
        x"31",
        x"50",
        x"54",
        x"53",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"51",
        x"45",
        x"42",
        x"09",
        x"0D",
        x"32",
        x"30",
        x"31",
        x"50",
        x"54",
        x"53",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"49",
        x"4D",
        x"42",
        x"09",
        x"0D",
        x"59",
        x"45",
        x"44",
        x"09",
        x"0D",
        x"59",
        x"45",
        x"44",
        x"09",
        x"0D",
        x"41",
        x"4D",
        x"41",
        x"4D",
        x"20",
        x"4F",
        x"4E",
        x"4F",
        x"53",
        x"09",
        x"09",
        x"30",
        x"31",
        x"31",
        x"50",
        x"54",
        x"53",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"51",
        x"45",
        x"42",
        x"09",
        x"0D",
        x"31",
        x"41",
        x"54",
        x"41",
        x"44",
        x"46",
        x"55",
        x"42",
        x"3A",
        x"20",
        x"5A",
        x"09",
        x"59",
        x"44",
        x"4C",
        x"09",
        x"31",
        x"53",
        x"50",
        x"4B",
        x"4E",
        x"54",
        x"53",
        x"0D",
        x"48",
        x"43",
        x"52",
        x"41",
        x"45",
        x"53",
        x"20",
        x"4B",
        x"4E",
        x"41",
        x"60",
        x"FF",
        x"49",
        x"0C",
        x"18",
        x"AD",
        x"0D",
        x"80",
        x"80",
        x"80",
        x"80",
        x"13",
        x"17",
        x"15",
        x"4F",
        x"11",
        x"80",
        x"80",
        x"10",
        x"4E",
        x"80",
        x"80",
        x"80",
        x"0C",
        x"0B",
        x"14",
        x"80",
        x"16",
        x"80",
        x"80",
        x"80",
        x"80",
        x"19",
        x"80",
        x"80",
        x"08",
        x"07",
        x"80",
        x"80",
        x"80",
        x"80",
        x"80",
        x"80",
        x"09",
        x"06",
        x"60",
        x"CE",
        x"D0",
        x"C5",
        x"C9",
        x"88",
        x"A5",
        x"E8",
        x"88",
        x"E6",
        x"02",
        x"30",
        x"0A",
        x"7F",
        x"41",
        x"BD",
        x"88",
        x"85",
        x"88",
        x"91",
        x"00",
        x"A0",
        x"88",
        x"84",
        x"88",
        x"A5",
        x"89",
        x"85",
        x"08",
        x"09",
        x"03",
        x"29",
        x"4A",
        x"4A",
        x"4A",
        x"7F",
        x"41",
        x"BD",
        x"A8",
        x"1A",
        x"09",
        x"0A",
        x"0A",
        x"0A",
        x"0A",
        x"0A",
        x"1E",
        x"30",
        x"7F",
        x"41",
        x"BD",
        x"00",
        x"A2",
        x"88",
        x"85",
        x"A0",
        x"A9",
        x"E1",
        x"D0",
        x"10",
        x"E0",
        x"E8",
        x"3D",
        x"B0",
        x"57",
        x"C0",
        x"41",
        x"90",
        x"4F",
        x"C0",
        x"00",
        x"B4",
        x"E8",
        x"48",
        x"B0",
        x"5F",
        x"C0",
        x"4C",
        x"90",
        x"57",
        x"C0",
        x"C8",
        x"01",
        x"90",
        x"0A",
        x"E0",
        x"00",
        x"B4",
        x"00",
        x"A2",
        x"60",
        x"18",
        x"98",
        x"60",
        x"F6",
        x"D0",
        x"04",
        x"C0",
        x"C8",
        x"06",
        x"10",
        x"0C",
        x"00",
        x"B9",
        x"00",
        x"A0",
        x"60",
        x"00",
        x"F6",
        x"60",
        x"00",
        x"D6",
        x"03",
        x"B0",
        x"E8",
        x"01",
        x"30",
        x"6A",
        x"6A",
        x"0C",
        x"B0",
        x"7E",
        x"D7",
        x"20",
        x"AA",
        x"0E",
        x"29",
        x"08",
        x"00",
        x"AD",
        x"60",
        x"08",
        x"00",
        x"EE",
        x"08",
        x"00",
        x"EE",
        x"06",
        x"D0",
        x"0C",
        x"C9",
        x"0F",
        x"29",
        x"08",
        x"01",
        x"8D",
        x"2A",
        x"08",
        x"01",
        x"AD",
        x"0A",
        x"0C",
        x"07",
        x"AD",
        x"7E",
        x"E7",
        x"20",
        x"7E",
        x"BF",
        x"20",
        x"7D",
        x"43",
        x"4C",
        x"F8",
        x"10",
        x"0C",
        x"0F",
        x"AD",
        x"0C",
        x"18",
        x"8D",
        x"68",
        x"66",
        x"4C",
        x"0E",
        x"85",
        x"B7",
        x"A9",
        x"0C",
        x"85",
        x"A7",
        x"A9",
        x"0A",
        x"85",
        x"97",
        x"A9",
        x"08",
        x"85",
        x"88",
        x"A9",
        x"06",
        x"85",
        x"78",
        x"A9",
        x"04",
        x"85",
        x"68",
        x"A9",
        x"02",
        x"85",
        x"58",
        x"A9",
        x"00",
        x"85",
        x"48",
        x"A9",
        x"0F",
        x"85",
        x"0D",
        x"85",
        x"0B",
        x"85",
        x"09",
        x"85",
        x"07",
        x"85",
        x"05",
        x"85",
        x"03",
        x"85",
        x"01",
        x"85",
        x"80",
        x"A9",
        x"35",
        x"D0",
        x"BF",
        x"C9",
        x"0A",
        x"02",
        x"AD",
        x"0A",
        x"E2",
        x"8D",
        x"C2",
        x"A9",
        x"0A",
        x"C2",
        x"8D",
        x"BF",
        x"A9",
        x"0A",
        x"A2",
        x"8D",
        x"BD",
        x"A9",
        x"0A",
        x"02",
        x"8D",
        x"A1",
        x"69",
        x"18",
        x"98",
        x"09",
        x"E2",
        x"8D",
        x"B0",
        x"A9",
        x"7E",
        x"48",
        x"4C",
        x"BF",
        x"A9",
        x"09",
        x"E2",
        x"8D",
        x"BB",
        x"A9",
        x"D6",
        x"D0",
        x"03",
        x"C0",
        x"0E",
        x"D0",
        x"7F",
        x"F5",
        x"D9",
        x"8A",
        x"A8",
        x"4A",
        x"4A",
        x"4A",
        x"60",
        x"E9",
        x"18",
        x"01",
        x"A5",
        x"ED",
        x"D0",
        x"07",
        x"29",
        x"01",
        x"A5",
        x"01",
        x"E6",
        x"AA",
        x"FA",
        x"D0",
        x"C8",
        x"00",
        x"71",
        x"18",
        x"8A",
        x"0C",
        x"18",
        x"8D",
        x"00",
        x"A0",
        x"00",
        x"A2",
        x"01",
        x"85",
        x"60",
        x"A9",
        x"00",
        x"85",
        x"00",
        x"A9",
        x"7D",
        x"43",
        x"4C",
        x"F8",
        x"10",
        x"0C",
        x"0F",
        x"AD",
        x"0C",
        x"18",
        x"8D",
        x"0B",
        x"F0",
        x"BF",
        x"C9",
        x"01",
        x"A5",
        x"0A",
        x"E4",
        x"8D",
        x"C2",
        x"A9",
        x"0A",
        x"C4",
        x"8D",
        x"B1",
        x"A9",
        x"0A",
        x"A4",
        x"8D",
        x"BD",
        x"A9",
        x"0A",
        x"04",
        x"8D",
        x"01",
        x"A5",
        x"09",
        x"E4",
        x"8D",
        x"00",
        x"A5",
        x"EE",
        x"D0",
        x"0C",
        x"C9",
        x"03",
        x"A5",
        x"03",
        x"E6",
        x"FB",
        x"D0",
        x"C8",
        x"02",
        x"91",
        x"0C",
        x"18",
        x"8D",
        x"B0",
        x"A9",
        x"A8",
        x"02",
        x"85",
        x"00",
        x"A9",
        x"03",
        x"85",
        x"08",
        x"A9",
        x"01",
        x"85",
        x"A1",
        x"69",
        x"18",
        x"4A",
        x"4A",
        x"01",
        x"A5",
        x"00",
        x"86",
        x"B8",
        x"A2",
        x"02",
        x"D0",
        x"0F",
        x"29",
        x"BC",
        x"A2",
        x"00",
        x"51",
        x"7D",
        x"BE",
        x"4C",
        x"01",
        x"85",
        x"BF",
        x"A9",
        x"00",
        x"85",
        x"BB",
        x"A9",
        x"BB",
        x"D0",
        x"10",
        x"E0",
        x"E8",
        x"02",
        x"A6",
        x"E8",
        x"D0",
        x"0C",
        x"C9",
        x"01",
        x"A5",
        x"01",
        x"E6",
        x"E8",
        x"AA",
        x"F6",
        x"D0",
        x"C8",
        x"11",
        x"69",
        x"18",
        x"22",
        x"D0",
        x"00",
        x"D1",
        x"8A",
        x"0C",
        x"18",
        x"8D",
        x"02",
        x"A6",
        x"02",
        x"A0",
        x"01",
        x"85",
        x"00",
        x"A9",
        x"EA",
        x"D0",
        x"0C",
        x"C9",
        x"01",
        x"A5",
        x"01",
        x"E6",
        x"E8",
        x"AA",
        x"F8",
        x"D0",
        x"C8",
        x"11",
        x"69",
        x"18",
        x"00",
        x"91",
        x"8A",
        x"0C",
        x"18",
        x"8D",
        x"02",
        x"A0",
        x"01",
        x"85",
        x"00",
        x"85",
        x"00",
        x"A9",
        x"00",
        x"A2",
        x"0C",
        x"0A",
        x"8C",
        x"C8",
        x"FB",
        x"D0",
        x"C8",
        x"00",
        x"91",
        x"A8",
        x"00",
        x"85",
        x"00",
        x"A9",
        x"01",
        x"85",
        x"D8",
        x"0C",
        x"A9",
        x"78",
        x"60",
        x"18",
        x"02",
        x"0B",
        x"AC",
        x"73",
        x"9A",
        x"20",
        x"60",
        x"A2",
        x"7A",
        x"A0",
        x"02",
        x"0B",
        x"8C",
        x"C2",
        x"D0",
        x"1A",
        x"C9",
        x"02",
        x"0A",
        x"AD",
        x"C9",
        x"D0",
        x"00",
        x"C9",
        x"02",
        x"09",
        x"AD",
        x"D0",
        x"D0",
        x"0F",
        x"C9",
        x"0F",
        x"29",
        x"02",
        x"08",
        x"AD",
        x"F2",
        x"D0",
        x"02",
        x"0B",
        x"CE",
        x"FA",
        x"10",
        x"CA",
        x"02",
        x"08",
        x"3E",
        x"4A",
        x"02",
        x"A2",
        x"02",
        x"0B",
        x"8E",
        x"02",
        x"A2",
        x"98",
        x"02",
        x"0F",
        x"8D",
        x"80",
        x"A9",
        x"F2",
        x"30",
        x"02",
        x"0F",
        x"2C",
        x"F7",
        x"30",
        x"0C",
        x"07",
        x"2C",
        x"F1",
        x"B0",
        x"60",
        x"18",
        x"60",
        x"02",
        x"0F",
        x"8D",
        x"00",
        x"A9",
        x"38",
        x"06",
        x"B0",
        x"04",
        x"E0",
        x"E0",
        x"D0",
        x"DB",
        x"F0",
        x"02",
        x"C9",
        x"C1",
        x"A5",
        x"40",
        x"0C",
        x"10",
        x"8D",
        x"68",
        x"AA",
        x"68",
        x"0C",
        x"02",
        x"8E",
        x"01",
        x"A2",
        x"02",
        x"B0",
        x"98",
        x"C9",
        x"C0",
        x"A5",
        x"00",
        x"A2",
        x"C8",
        x"85",
        x"30",
        x"A9",
        x"7B",
        x"A4",
        x"20",
        x"C1",
        x"85",
        x"00",
        x"A9",
        x"7B",
        x"A4",
        x"20",
        x"03",
        x"70",
        x"24",
        x"10",
        x"CB",
        x"24",
        x"C1",
        x"E6",
        x"0C",
        x"03",
        x"8D",
        x"70",
        x"B4",
        x"20",
        x"0C",
        x"03",
        x"8D",
        x"14",
        x"30",
        x"C6",
        x"24",
        x"20",
        x"A2",
        x"0C",
        x"08",
        x"8D",
        x"01",
        x"A9",
        x"EE",
        x"10",
        x"0C",
        x"07",
        x"AD",
        x"F3",
        x"10",
        x"0C",
        x"06",
        x"AD",
        x"F8",
        x"10",
        x"0C",
        x"05",
        x"AD",
        x"70",
        x"B4",
        x"20",
        x"C6",
        x"85",
        x"80",
        x"A9",
        x"40",
        x"30",
        x"0C",
        x"07",
        x"2C",
        x"07",
        x"10",
        x"0C",
        x"06",
        x"2C",
        x"0C",
        x"10",
        x"0C",
        x"05",
        x"2C",
        x"00",
        x"A9",
        x"0C",
        x"08",
        x"8E",
        x"03",
        x"D0",
        x"C8",
        x"86",
        x"CA",
        x"08",
        x"F0",
        x"C8",
        x"A6",
        x"0C",
        x"18",
        x"8D",
        x"48",
        x"8A",
        x"48",
        x"60",
        x"2A",
        x"91",
        x"00",
        x"A0",
        x"A0",
        x"09",
        x"2B",
        x"86",
        x"2A",
        x"84",
        x"DB",
        x"D0",
        x"60",
        x"A2",
        x"2C",
        x"A0",
        x"E1",
        x"D0",
        x"60",
        x"A2",
        x"38",
        x"A0",
        x"06",
        x"70",
        x"CB",
        x"24",
        x"73",
        x"9A",
        x"20",
        x"60",
        x"A2",
        x"14",
        x"A0",
        x"07",
        x"F0",
        x"73",
        x"9A",
        x"20",
        x"60",
        x"A2",
        x"20",
        x"A0",
        x"09",
        x"30",
        x"73",
        x"9A",
        x"4C",
        x"60",
        x"A2",
        x"44",
        x"A0",
        x"07",
        x"D0",
        x"CB",
        x"85",
        x"C0",
        x"29",
        x"6A",
        x"0C",
        x"19",
        x"0E",
        x"6A",
        x"0C",
        x"1A",
        x"0E",
        x"73",
        x"9A",
        x"20",
        x"60",
        x"A2",
        x"0A",
        x"A0",
        x"04",
        x"D0",
        x"60",
        x"A2",
        x"00",
        x"A0",
        x"06",
        x"10",
        x"CD",
        x"85",
        x"7F",
        x"68",
        x"20",
        x"73",
        x"9A",
        x"20",
        x"60",
        x"A2",
        x"69",
        x"A0",
        x"07",
        x"F0",
        x"6E",
        x"78",
        x"20",
        x"AA",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"60",
        x"A2",
        x"61",
        x"A0",
        x"0E",
        x"30",
        x"CC",
        x"A5",
        x"73",
        x"9A",
        x"20",
        x"60",
        x"A2",
        x"59",
        x"A0",
        x"CC",
        x"84",
        x"FF",
        x"A0",
        x"02",
        x"10",
        x"0C",
        x"1C",
        x"2C",
        x"20",
        x"A0",
        x"09",
        x"D0",
        x"15",
        x"A0",
        x"0D",
        x"10",
        x"0C",
        x"1C",
        x"2C",
        x"09",
        x"30",
        x"0C",
        x"1B",
        x"AD",
        x"10",
        x"A0",
        x"7C",
        x"61",
        x"20",
        x"09",
        x"A2",
        x"CC",
        x"A0",
        x"CA",
        x"85",
        x"03",
        x"A9",
        x"02",
        x"30",
        x"0C",
        x"1D",
        x"2C",
        x"02",
        x"A9",
        x"73",
        x"9A",
        x"20",
        x"60",
        x"A2",
        x"73",
        x"A0",
        x"CF",
        x"85",
        x"0C",
        x"1F",
        x"AD",
        x"CE",
        x"85",
        x"0C",
        x"1E",
        x"AD",
        x"60",
        x"D8",
        x"C0",
        x"85",
        x"01",
        x"E9",
        x"C0",
        x"A5",
        x"38",
        x"F8",
        x"60",
        x"D8",
        x"A0",
        x"95",
        x"A0",
        x"75",
        x"01",
        x"A9",
        x"18",
        x"F8",
        x"40",
        x"68",
        x"A8",
        x"68",
        x"AA",
        x"68",
        x"78",
        x"02",
        x"20",
        x"18",
        x"85",
        x"00",
        x"A9",
        x"17",
        x"85",
        x"06",
        x"49",
        x"8A",
        x"16",
        x"86",
        x"0E",
        x"F0",
        x"31",
        x"B5",
        x"04",
        x"A2",
        x"2C",
        x"02",
        x"A2",
        x"03",
        x"F0",
        x"02",
        x"29",
        x"8B",
        x"A5",
        x"7B",
        x"9E",
        x"4C",
        x"37",
        x"E6",
        x"78",
        x"02",
        x"20",
        x"18",
        x"85",
        x"0A",
        x"17",
        x"85",
        x"02",
        x"A9",
        x"16",
        x"86",
        x"00",
        x"A2",
        x"7B",
        x"9E",
        x"4C",
        x"12",
        x"46",
        x"02",
        x"F0",
        x"77",
        x"6F",
        x"20",
        x"3A",
        x"D0",
        x"76",
        x"5A",
        x"20",
        x"75",
        x"E5",
        x"20",
        x"0C",
        x"0C",
        x"8D",
        x"5A",
        x"85",
        x"11",
        x"A9",
        x"07",
        x"F0",
        x"B8",
        x"A5",
        x"37",
        x"86",
        x"00",
        x"A2",
        x"36",
        x"85",
        x"6C",
        x"A5",
        x"30",
        x"85",
        x"6D",
        x"A5",
        x"31",
        x"85",
        x"5B",
        x"F0",
        x"6E",
        x"A5",
        x"12",
        x"66",
        x"38",
        x"62",
        x"D0",
        x"77",
        x"6F",
        x"20",
        x"2D",
        x"30",
        x"12",
        x"24",
        x"3B",
        x"D0",
        x"31",
        x"A5",
        x"52",
        x"F0",
        x"01",
        x"29",
        x"8B",
        x"A5",
        x"75",
        x"10",
        x"8A",
        x"C6",
        x"04",
        x"F0",
        x"8A",
        x"A5",
        x"8F",
        x"85",
        x"00",
        x"A9",
        x"76",
        x"5A",
        x"20",
        x"75",
        x"E5",
        x"20",
        x"AA",
        x"98",
        x"31",
        x"96",
        x"AA",
        x"6E",
        x"B5",
        x"16",
        x"A6",
        x"30",
        x"96",
        x"AA",
        x"6D",
        x"B5",
        x"16",
        x"A6",
        x"36",
        x"96",
        x"AA",
        x"6C",
        x"B5",
        x"16",
        x"A6",
        x"02",
        x"A0",
        x"2C",
        x"04",
        x"A0",
        x"26",
        x"D0",
        x"35",
        x"A5",
        x"07",
        x"F0",
        x"33",
        x"A5",
        x"2E",
        x"B0",
        x"75",
        x"16",
        x"20",
        x"33",
        x"D0",
        x"8A",
        x"A4",
        x"37",
        x"10",
        x"58",
        x"24",
        x"04",
        x"B0",
        x"06",
        x"C0",
        x"04",
        x"30",
        x"CF",
        x"24",
        x"0C",
        x"B0",
        x"12",
        x"C0",
        x"68",
        x"A8",
        x"71",
        x"16",
        x"20",
        x"48",
        x"72",
        x"53",
        x"20",
        x"72",
        x"66",
        x"20",
        x"18",
        x"84",
        x"50",
        x"A0",
        x"16",
        x"A6",
        x"78",
        x"CF",
        x"20",
        x"1B",
        x"84",
        x"6D",
        x"A4",
        x"1C",
        x"84",
        x"06",
        x"D0",
        x"1C",
        x"84",
        x"6B",
        x"A4",
        x"1B",
        x"84",
        x"6A",
        x"A4",
        x"0A",
        x"F0",
        x"01",
        x"29",
        x"8A",
        x"05",
        x"F0",
        x"78",
        x"BC",
        x"20",
        x"76",
        x"D0",
        x"08",
        x"29",
        x"8B",
        x"A5",
        x"A7",
        x"D0",
        x"50",
        x"A0",
        x"16",
        x"A6",
        x"1D",
        x"85",
        x"66",
        x"B5",
        x"E8",
        x"01",
        x"F0",
        x"01",
        x"29",
        x"70",
        x"5E",
        x"20",
        x"1E",
        x"85",
        x"7B",
        x"A9",
        x"02",
        x"10",
        x"B5",
        x"24",
        x"63",
        x"A9",
        x"1F",
        x"85",
        x"63",
        x"B5",
        x"8E",
        x"85",
        x"57",
        x"85",
        x"00",
        x"A9",
        x"A5",
        x"E6",
        x"A6",
        x"E6",
        x"D9",
        x"D0",
        x"62",
        x"A1",
        x"AA",
        x"02",
        x"49",
        x"8A",
        x"08",
        x"F0",
        x"62",
        x"A1",
        x"AA",
        x"0A",
        x"01",
        x"29",
        x"70",
        x"5E",
        x"20",
        x"EC",
        x"10",
        x"57",
        x"24",
        x"41",
        x"D0",
        x"6E",
        x"B5",
        x"16",
        x"85",
        x"AA",
        x"1D",
        x"65",
        x"18",
        x"0A",
        x"1D",
        x"85",
        x"7B",
        x"21",
        x"4C",
        x"72",
        x"53",
        x"20",
        x"72",
        x"66",
        x"20",
        x"18",
        x"84",
        x"40",
        x"A0",
        x"00",
        x"A2",
        x"6D",
        x"91",
        x"C8",
        x"6D",
        x"91",
        x"20",
        x"A0",
        x"6D",
        x"91",
        x"C8",
        x"6D",
        x"91",
        x"A8",
        x"00",
        x"A9",
        x"0C",
        x"0B",
        x"8D",
        x"01",
        x"A9",
        x"5B",
        x"85",
        x"04",
        x"A9",
        x"06",
        x"F0",
        x"00",
        x"A9",
        x"0D",
        x"10",
        x"5B",
        x"C6",
        x"04",
        x"F0",
        x"5B",
        x"A5",
        x"1F",
        x"85",
        x"1E",
        x"86",
        x"1D",
        x"84",
        x"6E",
        x"A5",
        x"6D",
        x"A6",
        x"6C",
        x"A4",
        x"18",
        x"90",
        x"74",
        x"BA",
        x"20",
        x"6D",
        x"A4",
        x"6E",
        x"A6",
        x"98",
        x"0C",
        x"D0",
        x"6C",
        x"C4",
        x"0E",
        x"F0",
        x"6C",
        x"C4",
        x"12",
        x"30",
        x"5E",
        x"85",
        x"5E",
        x"A4",
        x"FF",
        x"A9",
        x"0C",
        x"90",
        x"79",
        x"A2",
        x"20",
        x"CF",
        x"F0",
        x"B8",
        x"A5",
        x"5F",
        x"F0",
        x"6E",
        x"A5",
        x"66",
        x"D0",
        x"07",
        x"29",
        x"8B",
        x"A5",
        x"5E",
        x"84",
        x"02",
        x"B0",
        x"79",
        x"A2",
        x"20",
        x"8B",
        x"E6",
        x"8D",
        x"E6",
        x"48",
        x"8A",
        x"48",
        x"98",
        x"48",
        x"7A",
        x"48",
        x"4C",
        x"78",
        x"CF",
        x"20",
        x"1C",
        x"85",
        x"09",
        x"A9",
        x"1B",
        x"85",
        x"E3",
        x"A9",
        x"78",
        x"BC",
        x"20",
        x"00",
        x"A2",
        x"01",
        x"03",
        x"00",
        x"02",
        x"FF",
        x"FF",
        x"FF",
        x"FF",
        x"00",
        x"02",
        x"01",
        x"03",
        x"60",
        x"A8",
        x"79",
        x"BC",
        x"BD",
        x"60",
        x"F6",
        x"10",
        x"88",
        x"04",
        x"90",
        x"0A",
        x"0C",
        x"00",
        x"BD",
        x"CA",
        x"0C",
        x"A2",
        x"02",
        x"10",
        x"B5",
        x"24",
        x"04",
        x"A2",
        x"03",
        x"A0",
        x"60",
        x"21",
        x"91",
        x"C8",
        x"21",
        x"91",
        x"20",
        x"A0",
        x"21",
        x"91",
        x"C8",
        x"21",
        x"91",
        x"A8",
        x"0A",
        x"58",
        x"85",
        x"00",
        x"A9",
        x"2C",
        x"80",
        x"A9",
        x"1F",
        x"86",
        x"1E",
        x"84",
        x"1D",
        x"85",
        x"21",
        x"A4",
        x"22",
        x"A6",
        x"20",
        x"A5",
        x"0F",
        x"90",
        x"74",
        x"BA",
        x"20",
        x"21",
        x"A4",
        x"22",
        x"A6",
        x"01",
        x"49",
        x"20",
        x"A5",
        x"1C",
        x"90",
        x"74",
        x"BA",
        x"20",
        x"21",
        x"A4",
        x"22",
        x"A6",
        x"01",
        x"49",
        x"1D",
        x"A5",
        x"29",
        x"90",
        x"74",
        x"BA",
        x"20",
        x"21",
        x"A4",
        x"22",
        x"A6",
        x"02",
        x"49",
        x"2C",
        x"03",
        x"49",
        x"03",
        x"30",
        x"28",
        x"20",
        x"A5",
        x"08",
        x"70",
        x"54",
        x"20",
        x"40",
        x"90",
        x"E6",
        x"B0",
        x"9B",
        x"C5",
        x"70",
        x"5E",
        x"20",
        x"46",
        x"90",
        x"0B",
        x"B0",
        x"9E",
        x"C5",
        x"61",
        x"A5",
        x"11",
        x"B0",
        x"74",
        x"BA",
        x"20",
        x"21",
        x"A4",
        x"22",
        x"A6",
        x"20",
        x"A5",
        x"13",
        x"90",
        x"74",
        x"BA",
        x"20",
        x"21",
        x"A4",
        x"22",
        x"A6",
        x"09",
        x"F0",
        x"20",
        x"C5",
        x"0D",
        x"30",
        x"17",
        x"B5",
        x"AA",
        x"01",
        x"49",
        x"8A",
        x"28",
        x"90",
        x"74",
        x"BE",
        x"20",
        x"1A",
        x"F0",
        x"20",
        x"C5",
        x"09",
        x"30",
        x"17",
        x"B5",
        x"AA",
        x"01",
        x"29",
        x"70",
        x"54",
        x"20",
        x"18",
        x"86",
        x"03",
        x"A2",
        x"2C",
        x"02",
        x"A2",
        x"03",
        x"B0",
        x"07",
        x"F0",
        x"18",
        x"C5",
        x"1F",
        x"29",
        x"21",
        x"A5",
        x"18",
        x"85",
        x"1F",
        x"29",
        x"1B",
        x"A5",
        x"80",
        x"A2",
        x"17",
        x"86",
        x"00",
        x"A2",
        x"2C",
        x"01",
        x"A2",
        x"03",
        x"B0",
        x"07",
        x"F0",
        x"17",
        x"C5",
        x"E0",
        x"29",
        x"21",
        x"A5",
        x"17",
        x"85",
        x"E0",
        x"29",
        x"1B",
        x"A5",
        x"80",
        x"A2",
        x"12",
        x"90",
        x"17",
        x"B0",
        x"04",
        x"F0",
        x"1C",
        x"C5",
        x"22",
        x"A5",
        x"60",
        x"22",
        x"84",
        x"1F",
        x"84",
        x"6E",
        x"B4",
        x"21",
        x"85",
        x"1E",
        x"85",
        x"6D",
        x"B5",
        x"20",
        x"85",
        x"1D",
        x"85",
        x"6C",
        x"B5",
        x"C8",
        x"10",
        x"19",
        x"B4",
        x"21",
        x"A6",
        x"00",
        x"A9",
        x"02",
        x"10",
        x"76",
        x"B0",
        x"20",
        x"21",
        x"86",
        x"78",
        x"41",
        x"4C",
        x"03",
        x"B0",
        x"76",
        x"DD",
        x"20",
        x"DD",
        x"10",
        x"FF",
        x"49",
        x"02",
        x"10",
        x"21",
        x"A5",
        x"1E",
        x"91",
        x"00",
        x"A0",
        x"FF",
        x"49",
        x"02",
        x"10",
        x"98",
        x"CB",
        x"D0",
        x"47",
        x"95",
        x"80",
        x"A9",
        x"77",
        x"90",
        x"20",
        x"D4",
        x"30",
        x"77",
        x"64",
        x"20",
        x"1E",
        x"91",
        x"1A",
        x"A4",
        x"98",
        x"1E",
        x"91",
        x"A8",
        x"00",
        x"A9",
        x"18",
        x"10",
        x"21",
        x"A5",
        x"1C",
        x"10",
        x"A8",
        x"30",
        x"B0",
        x"76",
        x"B0",
        x"20",
        x"00",
        x"A2",
        x"21",
        x"85",
        x"39",
        x"B0",
        x"76",
        x"B0",
        x"20",
        x"01",
        x"A2",
        x"60",
        x"76",
        x"4F",
        x"20",
        x"16",
        x"A6",
        x"9E",
        x"D0",
        x"19",
        x"A5",
        x"76",
        x"46",
        x"20",
        x"18",
        x"A6",
        x"00",
        x"B4",
        x"01",
        x"B5",
        x"16",
        x"A6",
        x"76",
        x"46",
        x"20",
        x"17",
        x"A6",
        x"00",
        x"B4",
        x"01",
        x"B5",
        x"16",
        x"A6",
        x"19",
        x"85",
        x"FF",
        x"A9",
        x"F1",
        x"10",
        x"CA",
        x"21",
        x"90",
        x"40",
        x"C9",
        x"2B",
        x"90",
        x"10",
        x"C9",
        x"08",
        x"F0",
        x"1B",
        x"B5",
        x"01",
        x"A2",
        x"B5",
        x"F0",
        x"80",
        x"E0",
        x"B9",
        x"F0",
        x"90",
        x"E0",
        x"08",
        x"B0",
        x"A0",
        x"C9",
        x"91",
        x"F0",
        x"50",
        x"C9",
        x"04",
        x"D0",
        x"50",
        x"E0",
        x"99",
        x"F0",
        x"0A",
        x"D0",
        x"40",
        x"C9",
        x"0E",
        x"D0",
        x"40",
        x"E0",
        x"0A",
        x"F0",
        x"16",
        x"A4",
        x"F0",
        x"29",
        x"35",
        x"F0",
        x"76",
        x"81",
        x"20",
        x"75",
        x"C5",
        x"20",
        x"16",
        x"A6",
        x"76",
        x"5F",
        x"4C",
        x"16",
        x"A6",
        x"62",
        x"D0",
        x"3C",
        x"95",
        x"6B",
        x"A5",
        x"3B",
        x"95",
        x"6A",
        x"A5",
        x"77",
        x"A9",
        x"20",
        x"13",
        x"85",
        x"48",
        x"95",
        x"C0",
        x"A9",
        x"75",
        x"30",
        x"77",
        x"64",
        x"20",
        x"7A",
        x"10",
        x"6E",
        x"95",
        x"19",
        x"A6",
        x"00",
        x"A9",
        x"77",
        x"A9",
        x"20",
        x"76",
        x"05",
        x"20",
        x"03",
        x"D0",
        x"13",
        x"85",
        x"13",
        x"05",
        x"48",
        x"95",
        x"58",
        x"A6",
        x"80",
        x"A9",
        x"0C",
        x"D0",
        x"19",
        x"A6",
        x"58",
        x"86",
        x"77",
        x"A0",
        x"20",
        x"26",
        x"30",
        x"77",
        x"37",
        x"20",
        x"78",
        x"41",
        x"4C",
        x"03",
        x"F0",
        x"77",
        x"06",
        x"20",
        x"60",
        x"0C",
        x"0D",
        x"8D",
        x"59",
        x"85",
        x"1F",
        x"A9",
        x"07",
        x"F0",
        x"B8",
        x"A5",
        x"60",
        x"3C",
        x"95",
        x"1F",
        x"A5",
        x"3B",
        x"95",
        x"1E",
        x"A5",
        x"74",
        x"96",
        x"20",
        x"03",
        x"D0",
        x"02",
        x"C0",
        x"74",
        x"AE",
        x"20",
        x"03",
        x"D0",
        x"01",
        x"C0",
        x"1D",
        x"A4",
        x"60",
        x"00",
        x"A9",
        x"02",
        x"90",
        x"D0",
        x"C9",
        x"70",
        x"5E",
        x"20",
        x"09",
        x"90",
        x"75",
        x"71",
        x"20",
        x"60",
        x"80",
        x"29",
        x"0C",
        x"04",
        x"BD",
        x"08",
        x"A2",
        x"02",
        x"10",
        x"B5",
        x"24",
        x"00",
        x"A2",
        x"0E",
        x"F0",
        x"B8",
        x"A5",
        x"60",
        x"F8",
        x"10",
        x"CA",
        x"CA",
        x"04",
        x"F0",
        x"3C",
        x"B5",
        x"0A",
        x"A2",
        x"19",
        x"86",
        x"ED",
        x"D0",
        x"1E",
        x"C5",
        x"6D",
        x"B5",
        x"F3",
        x"D0",
        x"1F",
        x"C5",
        x"F7",
        x"F0",
        x"6E",
        x"B5",
        x"1A",
        x"30",
        x"CA",
        x"CA",
        x"CA",
        x"18",
        x"A2",
        x"74",
        x"AE",
        x"20",
        x"77",
        x"4D",
        x"4C",
        x"74",
        x"96",
        x"20",
        x"74",
        x"AE",
        x"20",
        x"09",
        x"F0",
        x"05",
        x"30",
        x"88",
        x"88",
        x"12",
        x"F0",
        x"1B",
        x"A4",
        x"60",
        x"1C",
        x"C4",
        x"C8",
        x"C8",
        x"F5",
        x"D0",
        x"1B",
        x"C4",
        x"01",
        x"A0",
        x"06",
        x"F0",
        x"1B",
        x"C4",
        x"60",
        x"1C",
        x"C4",
        x"C8",
        x"03",
        x"D0",
        x"1B",
        x"C4",
        x"02",
        x"A0",
        x"06",
        x"F0",
        x"1B",
        x"C4",
        x"0E",
        x"D0",
        x"02",
        x"29",
        x"00",
        x"A0",
        x"1D",
        x"A5",
        x"1C",
        x"85",
        x"03",
        x"29",
        x"1C",
        x"A5",
        x"1B",
        x"85",
        x"03",
        x"29",
        x"1B",
        x"A5",
        x"60",
        x"38",
        x"60",
        x"18",
        x"F6",
        x"D0",
        x"20",
        x"C5",
        x"06",
        x"30",
        x"66",
        x"13",
        x"B9",
        x"88",
        x"20",
        x"85",
        x"1B",
        x"B5",
        x"AA",
        x"01",
        x"49",
        x"8A",
        x"A8",
        x"04",
        x"E9",
        x"38",
        x"03",
        x"F0",
        x"00",
        x"E0",
        x"10",
        x"A9",
        x"2C",
        x"08",
        x"A9",
        x"03",
        x"D0",
        x"02",
        x"29",
        x"1D",
        x"A5",
        x"60",
        x"18",
        x"FF",
        x"49",
        x"02",
        x"D0",
        x"65",
        x"CB",
        x"BE",
        x"65",
        x"EF",
        x"B9",
        x"A8",
        x"1B",
        x"75",
        x"18",
        x"FF",
        x"A9",
        x"2C",
        x"08",
        x"A9",
        x"2C",
        x"11",
        x"A9",
        x"2C",
        x"1A",
        x"A9",
        x"03",
        x"F0",
        x"08",
        x"30",
        x"88",
        x"88",
        x"0F",
        x"F0",
        x"1D",
        x"A4",
        x"F7",
        x"B0",
        x"10",
        x"C9",
        x"FA",
        x"F0",
        x"1B",
        x"B5",
        x"60",
        x"38",
        x"60",
        x"1C",
        x"05",
        x"98",
        x"AA",
        x"F0",
        x"29",
        x"1C",
        x"25",
        x"A8",
        x"1B",
        x"85",
        x"1E",
        x"B1",
        x"19",
        x"84",
        x"00",
        x"A0",
        x"1C",
        x"85",
        x"1A",
        x"84",
        x"1E",
        x"B1",
        x"20",
        x"A0",
        x"2C",
        x"01",
        x"A0",
        x"03",
        x"D0",
        x"02",
        x"29",
        x"1D",
        x"85",
        x"36",
        x"B5",
        x"1F",
        x"85",
        x"31",
        x"B5",
        x"1E",
        x"85",
        x"30",
        x"B5",
        x"60",
        x"00",
        x"95",
        x"00",
        x"75",
        x"18",
        x"19",
        x"A5",
        x"60",
        x"00",
        x"95",
        x"1A",
        x"E5",
        x"38",
        x"00",
        x"B5",
        x"08",
        x"F0",
        x"01",
        x"29",
        x"E8",
        x"01",
        x"90",
        x"02",
        x"C9",
        x"36",
        x"B5",
        x"1A",
        x"84",
        x"19",
        x"85",
        x"A8",
        x"04",
        x"A9",
        x"03",
        x"D0",
        x"A8",
        x"08",
        x"A9",
        x"60",
        x"19",
        x"85",
        x"00",
        x"95",
        x"01",
        x"95",
        x"31",
        x"95",
        x"00",
        x"A9",
        x"0A",
        x"D0",
        x"00",
        x"D5",
        x"98",
        x"0F",
        x"D0",
        x"01",
        x"D5",
        x"60",
        x"D8",
        x"54",
        x"85",
        x"00",
        x"69",
        x"54",
        x"A5",
        x"53",
        x"85",
        x"53",
        x"65",
        x"18",
        x"F8",
        x"0D",
        x"F0",
        x"B8",
        x"A4",
        x"F7",
        x"D0",
        x"0A",
        x"A9",
        x"60",
        x"48",
        x"95",
        x"58",
        x"A6",
        x"05",
        x"F0",
        x"0C",
        x"C0",
        x"09",
        x"F0",
        x"06",
        x"C0",
        x"A7",
        x"A4",
        x"0A",
        x"D0",
        x"08",
        x"C9",
        x"02",
        x"69",
        x"10",
        x"D0",
        x"28",
        x"06",
        x"49",
        x"06",
        x"29",
        x"4A",
        x"4A",
        x"4A",
        x"0B",
        x"69",
        x"37",
        x"A5",
        x"08",
        x"18",
        x"1D",
        x"C5",
        x"01",
        x"49",
        x"6C",
        x"B5",
        x"60",
        x"01",
        x"95",
        x"06",
        x"69",
        x"18",
        x"0A",
        x"0A",
        x"0A",
        x"30",
        x"B5",
        x"00",
        x"95",
        x"01",
        x"E9",
        x"38",
        x"F8",
        x"49",
        x"F8",
        x"29",
        x"6A",
        x"1E",
        x"46",
        x"6A",
        x"1E",
        x"46",
        x"30",
        x"B5",
        x"1E",
        x"85",
        x"31",
        x"B5",
        x"60",
        x"30",
        x"95",
        x"1E",
        x"65",
        x"18",
        x"4A",
        x"4A",
        x"4A",
        x"01",
        x"B5",
        x"31",
        x"95",
        x"2A",
        x"1E",
        x"06",
        x"2A",
        x"1E",
        x"06",
        x"02",
        x"A9",
        x"1E",
        x"85",
        x"F8",
        x"29",
        x"F8",
        x"49",
        x"03",
        x"69",
        x"18",
        x"00",
        x"B5",
        x"60",
        x"01",
        x"A9",
        x"18",
        x"EF",
        x"10",
        x"CA",
        x"04",
        x"F0",
        x"50",
        x"C9",
        x"F0",
        x"29",
        x"F1",
        x"90",
        x"0B",
        x"F0",
        x"10",
        x"C9",
        x"1B",
        x"B5",
        x"01",
        x"A2",
        x"FB",
        x"F0",
        x"60",
        x"00",
        x"A9",
        x"60",
        x"F8",
        x"F0",
        x"75",
        x"AC",
        x"20",
        x"75",
        x"09",
        x"20",
        x"60",
        x"F8",
        x"F0",
        x"75",
        x"AC",
        x"20",
        x"75",
        x"01",
        x"20",
        x"60",
        x"F8",
        x"F0",
        x"75",
        x"AC",
        x"20",
        x"74",
        x"F5",
        x"20",
        x"60",
        x"F8",
        x"F0",
        x"75",
        x"AC",
        x"20",
        x"74",
        x"C9",
        x"20",
        x"1B",
        x"F0",
        x"14",
        x"30",
        x"88",
        x"88",
        x"0F",
        x"F0",
        x"1D",
        x"84",
        x"6C",
        x"A4",
        x"1F",
        x"84",
        x"6E",
        x"A4",
        x"1E",
        x"84",
        x"6D",
        x"A4",
        x"60",
        x"01",
        x"A9",
        x"9C",
        x"C5",
        x"60",
        x"A5",
        x"60",
        x"01",
        x"A9",
        x"8F",
        x"C5",
        x"9D",
        x"A5",
        x"E7",
        x"10",
        x"CA",
        x"0A",
        x"F0",
        x"40",
        x"C9",
        x"0E",
        x"F0",
        x"80",
        x"C9",
        x"12",
        x"F0",
        x"90",
        x"C9",
        x"F0",
        x"29",
        x"F1",
        x"90",
        x"13",
        x"F0",
        x"10",
        x"C9",
        x"1B",
        x"B5",
        x"01",
        x"A2",
        x"FB",
        x"F0",
        x"60",
        x"00",
        x"A9",
        x"60",
        x"F8",
        x"F0",
        x"75",
        x"46",
        x"20",
        x"75",
        x"09",
        x"20",
        x"60",
        x"F8",
        x"F0",
        x"75",
        x"46",
        x"20",
        x"75",
        x"01",
        x"20",
        x"60",
        x"F8",
        x"F0",
        x"75",
        x"46",
        x"20",
        x"74",
        x"F5",
        x"20",
        x"60",
        x"F8",
        x"F0",
        x"75",
        x"46",
        x"20",
        x"74",
        x"C9",
        x"20",
        x"1B",
        x"F0",
        x"14",
        x"30",
        x"88",
        x"88",
        x"0F",
        x"F0",
        x"A8",
        x"BE",
        x"D0",
        x"21",
        x"A0",
        x"1B",
        x"85",
        x"1E",
        x"B1",
        x"01",
        x"A0",
        x"74",
        x"86",
        x"20",
        x"74",
        x"FA",
        x"4C",
        x"74",
        x"A2",
        x"20",
        x"20",
        x"A0",
        x"D3",
        x"D0",
        x"C8",
        x"1B",
        x"85",
        x"1E",
        x"B1",
        x"74",
        x"AE",
        x"20",
        x"00",
        x"A0",
        x"60",
        x"AA",
        x"38",
        x"60",
        x"18",
        x"ED",
        x"10",
        x"CA",
        x"05",
        x"90",
        x"A0",
        x"C0",
        x"04",
        x"90",
        x"80",
        x"C0",
        x"0D",
        x"90",
        x"60",
        x"C0",
        x"0C",
        x"F0",
        x"1B",
        x"B4",
        x"01",
        x"A2",
        x"8A",
        x"1B",
        x"05",
        x"1C",
        x"85",
        x"1E",
        x"B1",
        x"20",
        x"A0",
        x"1B",
        x"85",
        x"1E",
        x"B1",
        x"74",
        x"96",
        x"20",
        x"00",
        x"A0",
        x"40",
        x"F0",
        x"3A",
        x"30",
        x"88",
        x"88",
        x"34",
        x"F0",
        x"A8",
        x"1D",
        x"85",
        x"1E",
        x"84",
        x"1F",
        x"86",
        x"60",
        x"1E",
        x"85",
        x"1F",
        x"C6",
        x"02",
        x"B0",
        x"20",
        x"E9",
        x"1E",
        x"A5",
        x"38",
        x"60",
        x"1E",
        x"85",
        x"1F",
        x"E6",
        x"02",
        x"90",
        x"20",
        x"69",
        x"1E",
        x"A5",
        x"18",
        x"60",
        x"1E",
        x"85",
        x"1F",
        x"C6",
        x"02",
        x"B0",
        x"01",
        x"E9",
        x"1E",
        x"A5",
        x"38",
        x"60",
        x"22",
        x"E6",
        x"02",
        x"D0",
        x"21",
        x"E6",
        x"21",
        x"91",
        x"60",
        x"1F",
        x"E6",
        x"02",
        x"D0",
        x"1E",
        x"E6",
        x"60",
        x"28",
        x"85",
        x"29",
        x"C6",
        x"02",
        x"B0",
        x"20",
        x"E9",
        x"28",
        x"A5",
        x"38",
        x"60",
        x"28",
        x"85",
        x"29",
        x"E6",
        x"02",
        x"90",
        x"20",
        x"69",
        x"28",
        x"A5",
        x"18",
        x"60",
        x"23",
        x"85",
        x"04",
        x"A9",
        x"AA",
        x"0A",
        x"0A",
        x"0A",
        x"8A",
        x"60",
        x"00",
        x"A9",
        x"02",
        x"B0",
        x"90",
        x"C9",
        x"06",
        x"90",
        x"11",
        x"C9",
        x"28",
        x"B1",
        x"E8",
        x"C8",
        x"60",
        x"10",
        x"A9",
        x"05",
        x"D0",
        x"1D",
        x"C9",
        x"04",
        x"F0",
        x"02",
        x"C9",
        x"1F",
        x"29",
        x"28",
        x"65",
        x"18",
        x"98",
        x"0E",
        x"90",
        x"5E",
        x"C9",
        x"28",
        x"A5",
        x"06",
        x"D0",
        x"08",
        x"C9",
        x"18",
        x"B0",
        x"0C",
        x"90",
        x"A2",
        x"C9",
        x"28",
        x"A5",
        x"08",
        x"D0",
        x"0B",
        x"C9",
        x"29",
        x"A5",
        x"60",
        x"28",
        x"91",
        x"01",
        x"69",
        x"C8",
        x"28",
        x"91",
        x"01",
        x"69",
        x"20",
        x"A0",
        x"28",
        x"91",
        x"01",
        x"69",
        x"C8",
        x"28",
        x"91",
        x"18",
        x"00",
        x"A0",
        x"2E",
        x"65",
        x"18",
        x"29",
        x"84",
        x"09",
        x"A0",
        x"28",
        x"84",
        x"FB",
        x"A0",
        x"80",
        x"A9",
        x"F6",
        x"30",
        x"B5",
        x"24",
        x"08",
        x"D0",
        x"E3",
        x"A0",
        x"90",
        x"A9",
        x"12",
        x"D0",
        x"2E",
        x"86",
        x"0C",
        x"A2",
        x"90",
        x"A9",
        x"09",
        x"A0",
        x"28",
        x"84",
        x"C0",
        x"A0",
        x"09",
        x"A1",
        x"8E",
        x"E8",
        x"09",
        x"A0",
        x"8E",
        x"9A",
        x"A2",
        x"11",
        x"D0",
        x"80",
        x"A9",
        x"0A",
        x"A0",
        x"28",
        x"84",
        x"1E",
        x"A0",
        x"0A",
        x"5F",
        x"8E",
        x"E8",
        x"0A",
        x"5E",
        x"8E",
        x"8A",
        x"A2",
        x"26",
        x"D0",
        x"0C",
        x"A0",
        x"80",
        x"A9",
        x"00",
        x"A2",
        x"60",
        x"29",
        x"85",
        x"3C",
        x"B5",
        x"28",
        x"85",
        x"3B",
        x"B5",
        x"60",
        x"F6",
        x"D0",
        x"88",
        x"74",
        x"7A",
        x"20",
        x"28",
        x"81",
        x"2A",
        x"B1",
        x"00",
        x"A2",
        x"A8",
        x"2A",
        x"B1",
        x"2B",
        x"E6",
        x"02",
        x"D0",
        x"2A",
        x"E6",
        x"29",
        x"85",
        x"2A",
        x"B1",
        x"2B",
        x"E6",
        x"02",
        x"D0",
        x"2A",
        x"E6",
        x"28",
        x"85",
        x"2A",
        x"B1",
        x"00",
        x"A0",
        x"2A",
        x"84",
        x"2B",
        x"86",
        x"60",
        x"E5",
        x"D0",
        x"23",
        x"C6",
        x"74",
        x"96",
        x"20",
        x"F2",
        x"D0",
        x"CA",
        x"74",
        x"8D",
        x"20",
        x"01",
        x"A9",
        x"02",
        x"90",
        x"00",
        x"A9",
        x"24",
        x"46",
        x"24",
        x"85",
        x"1E",
        x"B1",
        x"08",
        x"A2",
        x"04",
        x"10",
        x"4A",
        x"4A",
        x"4A",
        x"4A",
        x"1E",
        x"B1",
        x"04",
        x"A2",
        x"23",
        x"86",
        x"55",
        x"A2",
        x"00",
        x"A0",
        x"22",
        x"86",
        x"21",
        x"84",
        x"05",
        x"A2",
        x"40",
        x"A0",
        x"1F",
        x"85",
        x"1E",
        x"84",
        x"62",
        x"18",
        x"BD",
        x"A8",
        x"62",
        x"17",
        x"BD",
        x"72",
        x"EF",
        x"20",
        x"B4",
        x"10",
        x"CD",
        x"24",
        x"60",
        x"BA",
        x"86",
        x"E5",
        x"D0",
        x"23",
        x"C6",
        x"74",
        x"86",
        x"20",
        x"F2",
        x"D0",
        x"CA",
        x"74",
        x"8D",
        x"20",
        x"01",
        x"A9",
        x"02",
        x"90",
        x"00",
        x"A9",
        x"24",
        x"06",
        x"24",
        x"85",
        x"1E",
        x"B1",
        x"08",
        x"A2",
        x"23",
        x"86",
        x"55",
        x"A2",
        x"00",
        x"A0",
        x"22",
        x"86",
        x"21",
        x"84",
        x"05",
        x"A2",
        x"40",
        x"A0",
        x"04",
        x"F0",
        x"BA",
        x"A5",
        x"04",
        x"D0",
        x"B5",
        x"A5",
        x"02",
        x"A2",
        x"80",
        x"A0",
        x"1E",
        x"84",
        x"1F",
        x"85",
        x"62",
        x"08",
        x"BD",
        x"A8",
        x"62",
        x"07",
        x"BD",
        x"72",
        x"EF",
        x"20",
        x"BA",
        x"C6",
        x"60",
        x"AA",
        x"0A",
        x"61",
        x"FE",
        x"BD",
        x"03",
        x"30",
        x"CF",
        x"24",
        x"61",
        x"F5",
        x"BD",
        x"0A",
        x"10",
        x"07",
        x"29",
        x"C2",
        x"A5",
        x"06",
        x"90",
        x"09",
        x"E0",
        x"A3",
        x"A6",
        x"F7",
        x"F0",
        x"B8",
        x"A5",
        x"72",
        x"FB",
        x"4C",
        x"C7",
        x"A5",
        x"60",
        x"08",
        x"C9",
        x"1F",
        x"A5",
        x"04",
        x"D0",
        x"42",
        x"C9",
        x"74",
        x"AE",
        x"20",
        x"60",
        x"E8",
        x"D0",
        x"72",
        x"DE",
        x"20",
        x"F1",
        x"D0",
        x"24",
        x"C6",
        x"74",
        x"8F",
        x"20",
        x"1E",
        x"91",
        x"24",
        x"A4",
        x"21",
        x"B1",
        x"00",
        x"A0",
        x"24",
        x"84",
        x"1A",
        x"A0",
        x"72",
        x"81",
        x"20",
        x"05",
        x"A2",
        x"40",
        x"A0",
        x"04",
        x"D0",
        x"02",
        x"A2",
        x"80",
        x"A0",
        x"60",
        x"E4",
        x"D0",
        x"72",
        x"DE",
        x"20",
        x"ED",
        x"D0",
        x"24",
        x"C6",
        x"74",
        x"8D",
        x"20",
        x"00",
        x"A0",
        x"00",
        x"A9",
        x"02",
        x"90",
        x"11",
        x"C9",
        x"1E",
        x"B1",
        x"24",
        x"A4",
        x"24",
        x"84",
        x"1A",
        x"A0",
        x"72",
        x"81",
        x"20",
        x"05",
        x"A2",
        x"40",
        x"A0",
        x"04",
        x"D0",
        x"02",
        x"A2",
        x"80",
        x"A0",
        x"60",
        x"1F",
        x"86",
        x"1E",
        x"84",
        x"0B",
        x"A2",
        x"82",
        x"A0",
        x"22",
        x"86",
        x"21",
        x"84",
        x"60",
        x"1E",
        x"91",
        x"01",
        x"69",
        x"C8",
        x"1E",
        x"91",
        x"20",
        x"A0",
        x"01",
        x"69",
        x"1E",
        x"91",
        x"C8",
        x"01",
        x"69",
        x"1E",
        x"91",
        x"00",
        x"A0",
        x"18",
        x"65",
        x"0A",
        x"0A",
        x"1D",
        x"A5",
        x"1D",
        x"85",
        x"1E",
        x"84",
        x"1F",
        x"86",
        x"60",
        x"6C",
        x"95",
        x"1D",
        x"A5",
        x"6E",
        x"95",
        x"1F",
        x"A5",
        x"6D",
        x"95",
        x"1E",
        x"A5",
        x"60",
        x"A8",
        x"25",
        x"65",
        x"18",
        x"98",
        x"2A",
        x"91",
        x"00",
        x"A9",
        x"02",
        x"30",
        x"26",
        x"24",
        x"A0",
        x"09",
        x"2C",
        x"D0",
        x"09",
        x"03",
        x"10",
        x"B5",
        x"24",
        x"26",
        x"C6",
        x"02",
        x"F0",
        x"60",
        x"E5",
        x"10",
        x"2D",
        x"C6",
        x"CA",
        x"72",
        x"38",
        x"20",
        x"0F",
        x"29",
        x"68",
        x"26",
        x"C6",
        x"02",
        x"D0",
        x"2D",
        x"A5",
        x"72",
        x"38",
        x"20",
        x"4A",
        x"4A",
        x"4A",
        x"4A",
        x"48",
        x"A0",
        x"B5",
        x"26",
        x"85",
        x"00",
        x"A9",
        x"2D",
        x"85",
        x"02",
        x"A9",
        x"2A",
        x"85",
        x"A0",
        x"A0",
        x"25",
        x"84",
        x"E0",
        x"A0",
        x"2B",
        x"84",
        x"08",
        x"F0",
        x"00",
        x"A0",
        x"25",
        x"84",
        x"20",
        x"A0",
        x"2B",
        x"84",
        x"09",
        x"A0",
        x"9E",
        x"A9",
        x"25",
        x"A2",
        x"06",
        x"D0",
        x"08",
        x"A0",
        x"5E",
        x"A9",
        x"42",
        x"A2",
        x"0E",
        x"D0",
        x"0A",
        x"A0",
        x"BE",
        x"A9",
        x"5A",
        x"A2",
        x"20",
        x"D0",
        x"09",
        x"A0",
        x"C1",
        x"A9",
        x"25",
        x"A2",
        x"28",
        x"D0",
        x"0B",
        x"A0",
        x"01",
        x"A9",
        x"42",
        x"A2",
        x"30",
        x"D0",
        x"08",
        x"A0",
        x"A1",
        x"A9",
        x"5A",
        x"A2",
        x"28",
        x"30",
        x"71",
        x"F2",
        x"20",
        x"71",
        x"EA",
        x"20",
        x"0B",
        x"7E",
        x"8D",
        x"0B",
        x"5E",
        x"8D",
        x"09",
        x"1E",
        x"8D",
        x"08",
        x"FE",
        x"8D",
        x"0A",
        x"5E",
        x"8D",
        x"0A",
        x"3E",
        x"8D",
        x"D0",
        x"A9",
        x"2C",
        x"30",
        x"71",
        x"DA",
        x"20",
        x"71",
        x"D2",
        x"20",
        x"08",
        x"A1",
        x"8D",
        x"08",
        x"81",
        x"8D",
        x"09",
        x"D0",
        x"C9",
        x"A4",
        x"0B",
        x"01",
        x"8D",
        x"0A",
        x"E1",
        x"8D",
        x"09",
        x"C1",
        x"8D",
        x"09",
        x"A1",
        x"8D",
        x"A0",
        x"A9",
        x"60",
        x"AA",
        x"26",
        x"65",
        x"0A",
        x"0A",
        x"60",
        x"9B",
        x"85",
        x"65",
        x"8F",
        x"BD",
        x"71",
        x"90",
        x"20",
        x"95",
        x"A5",
        x"9E",
        x"85",
        x"65",
        x"BF",
        x"BD",
        x"71",
        x"90",
        x"20",
        x"98",
        x"A5",
        x"9D",
        x"85",
        x"65",
        x"AF",
        x"BD",
        x"71",
        x"90",
        x"20",
        x"97",
        x"A5",
        x"9C",
        x"85",
        x"65",
        x"9F",
        x"BD",
        x"71",
        x"90",
        x"20",
        x"96",
        x"A5",
        x"9A",
        x"85",
        x"65",
        x"7F",
        x"BD",
        x"71",
        x"90",
        x"20",
        x"94",
        x"A5",
        x"99",
        x"85",
        x"65",
        x"6F",
        x"BD",
        x"71",
        x"90",
        x"20",
        x"93",
        x"A5",
        x"A7",
        x"85",
        x"A6",
        x"85",
        x"A5",
        x"85",
        x"00",
        x"A9",
        x"F0",
        x"10",
        x"CA",
        x"C8",
        x"93",
        x"95",
        x"65",
        x"1F",
        x"B9",
        x"03",
        x"30",
        x"CF",
        x"24",
        x"64",
        x"CF",
        x"B9",
        x"05",
        x"A2",
        x"A8",
        x"0A",
        x"0A",
        x"0A",
        x"09",
        x"A9",
        x"02",
        x"90",
        x"0A",
        x"C9",
        x"71",
        x"16",
        x"20",
        x"26",
        x"85",
        x"6F",
        x"B5",
        x"20",
        x"7B",
        x"A4",
        x"20",
        x"03",
        x"A2",
        x"60",
        x"D8",
        x"03",
        x"69",
        x"18",
        x"F8",
        x"05",
        x"30",
        x"CE",
        x"24",
        x"A3",
        x"A5",
        x"60",
        x"68",
        x"F6",
        x"D0",
        x"CA",
        x"74",
        x"AE",
        x"20",
        x"48",
        x"1E",
        x"91",
        x"68",
        x"1B",
        x"A2",
        x"00",
        x"A0",
        x"1F",
        x"84",
        x"0B",
        x"A0",
        x"1E",
        x"84",
        x"48",
        x"9D",
        x"A0",
        x"70",
        x"FF",
        x"20",
        x"82",
        x"A0",
        x"70",
        x"DE",
        x"20",
        x"A2",
        x"A0",
        x"0B",
        x"A2",
        x"70",
        x"DC",
        x"20",
        x"42",
        x"A0",
        x"08",
        x"A2",
        x"60",
        x"FB",
        x"10",
        x"88",
        x"1E",
        x"91",
        x"1B",
        x"A0",
        x"1F",
        x"86",
        x"1E",
        x"84",
        x"10",
        x"A9",
        x"60",
        x"DC",
        x"D0",
        x"28",
        x"68",
        x"6C",
        x"1D",
        x"4C",
        x"03",
        x"F0",
        x"C0",
        x"A5",
        x"07",
        x"30",
        x"B8",
        x"A5",
        x"7D",
        x"43",
        x"4C",
        x"03",
        x"30",
        x"0C",
        x"0F",
        x"AD",
        x"48",
        x"08",
        x"0C",
        x"18",
        x"8D",
        x"01",
        x"E9",
        x"68",
        x"FC",
        x"D0",
        x"01",
        x"E9",
        x"48",
        x"38",
        x"50",
        x"A9",
        x"2C",
        x"0C",
        x"0D",
        x"8D",
        x"0C",
        x"0C",
        x"8D",
        x"0C",
        x"09",
        x"8D",
        x"00",
        x"A9",
        x"0C",
        x"0A",
        x"8D",
        x"01",
        x"A9",
        x"60",
        x"FA",
        x"D0",
        x"CA",
        x"70",
        x"A3",
        x"20",
        x"0D",
        x"A2",
        x"2C",
        x"06",
        x"A2",
        x"2C",
        x"04",
        x"A2",
        x"60",
        x"F6",
        x"D0",
        x"1F",
        x"A5",
        x"0C",
        x"18",
        x"8D",
        x"74",
        x"96",
        x"20",
        x"1F",
        x"85",
        x"C0",
        x"A9",
        x"2C",
        x"03",
        x"A9",
        x"60",
        x"C2",
        x"85",
        x"60",
        x"A5",
        x"61",
        x"85",
        x"61",
        x"65",
        x"43",
        x"A9",
        x"06",
        x"D0",
        x"60",
        x"25",
        x"4A",
        x"A9",
        x"60",
        x"66",
        x"61",
        x"66",
        x"4A",
        x"00",
        x"69",
        x"61",
        x"25",
        x"01",
        x"A9",
        x"38",
        x"01",
        x"F0",
        x"18",
        x"60",
        x"25",
        x"02",
        x"A9",
        x"60",
        x"FF",
        x"49",
        x"02",
        x"10",
        x"B5",
        x"24",
        x"70",
        x"5E",
        x"20",
        x"60",
        x"DB",
        x"90",
        x"C0",
        x"C9",
        x"28",
        x"A5",
        x"E1",
        x"D0",
        x"0B",
        x"C9",
        x"29",
        x"A5",
        x"74",
        x"6E",
        x"20",
        x"EC",
        x"90",
        x"1F",
        x"C0",
        x"74",
        x"24",
        x"20",
        x"18",
        x"DA",
        x"A9",
        x"2C",
        x"EA",
        x"A9",
        x"03",
        x"F0",
        x"20",
        x"29",
        x"28",
        x"A5",
        x"C8",
        x"FF",
        x"A0",
        x"29",
        x"86",
        x"28",
        x"84",
        x"08",
        x"A2",
        x"40",
        x"A0",
        x"60",
        x"F6",
        x"D0",
        x"CA",
        x"1F",
        x"C6",
        x"FB",
        x"D0",
        x"1E",
        x"91",
        x"88",
        x"04",
        x"A2",
        x"1E",
        x"84",
        x"00",
        x"A0",
        x"1F",
        x"84",
        x"0B",
        x"A0",
        x"00",
        x"A9",
        x"FB",
        x"10",
        x"CA",
        x"00",
        x"95",
        x"0F",
        x"A2",
        x"00",
        x"A9",
        x"60",
        x"F8",
        x"10",
        x"88",
        x"CA",
        x"60",
        x"95",
        x"1E",
        x"B1",
        x"23",
        x"A6",
        x"1E",
        x"85",
        x"1F",
        x"86",
        x"23",
        x"84",
        x"0E",
        x"A0",
        x"32",
        x"A9",
        x"66",
        x"A2",
        x"04",
        x"D0",
        x"23",
        x"A9",
        x"66",
        x"A2",
        x"EB",
        x"D0",
        x"23",
        x"84",
        x"47",
        x"A0",
        x"00",
        x"A2",
        x"E8",
        x"A9",
        x"2C",
        x"D0",
        x"A9",
        x"1B",
        x"D0",
        x"17",
        x"A0",
        x"2D",
        x"F0",
        x"B8",
        x"A4",
        x"90",
        x"A9",
        x"00",
        x"A2",
        x"23",
        x"85",
        x"9F",
        x"A9",
        x"2C",
        x"87",
        x"A9",
        x"60",
        x"0C",
        x"0A",
        x"8E",
        x"E8",
        x"0C",
        x"09",
        x"8E",
        x"F8",
        x"D0",
        x"0C",
        x"18",
        x"8D",
        x"00",
        x"95",
        x"CA",
        x"00",
        x"A9",
        x"9F",
        x"A2",
        x"2C",
        x"C0",
        x"A2",
        x"2C",
        x"00",
        x"A2",
        x"12",
        x"F0",
        x"F8",
        x"D0",
        x"0C",
        x"18",
        x"8D",
        x"10",
        x"95",
        x"CA",
        x"00",
        x"A9",
        x"F0",
        x"A2",
        x"60",
        x"FA",
        x"10",
        x"CA",
        x"0C",
        x"00",
        x"9D",
        x"00",
        x"A9",
        x"18",
        x"A2",
        x"60",
        x"0C",
        x"00",
        x"8E",
        x"0C",
        x"01",
        x"8E",
        x"E8",
        x"B8",
        x"86",
        x"FF",
        x"A2",
        x"7B",
        x"AE",
        x"20",
        x"7B",
        x"AE",
        x"20",
        x"03",
        x"50",
        x"08",
        x"F0",
        x"CB",
        x"A5",
        x"C9",
        x"84",
        x"B4",
        x"84",
        x"40",
        x"A0",
        x"02",
        x"70",
        x"00",
        x"A0",
        x"F0",
        x"90",
        x"02",
        x"F0",
        x"CB",
        x"A5",
        x"01",
        x"E0",
        x"AD",
        x"02",
        x"E0",
        x"BA",
        x"F0",
        x"E8",
        x"D0",
        x"88",
        x"05",
        x"10",
        x"0A",
        x"50",
        x"5F",
        x"24",
        x"5F",
        x"85",
        x"6A",
        x"0C",
        x"0E",
        x"0E",
        x"6A",
        x"0C",
        x"0D",
        x"0E",
        x"C0",
        x"A6",
        x"70",
        x"B4",
        x"20",
        x"10",
        x"A0",
        x"0C",
        x"00",
        x"8D",
        x"0C",
        x"01",
        x"8D",
        x"03",
        x"F0",
        x"01",
        x"E0",
        x"C0",
        x"A6",
        x"27",
        x"85",
        x"01",
        x"49",
        x"27",
        x"A5",
        x"6E",
        x"E8",
        x"20",
        x"7B",
        x"A4",
        x"20",
        x"03",
        x"A2",
        x"08",
        x"D0",
        x"77",
        x"73",
        x"20",
        x"0D",
        x"D0",
        x"CB",
        x"A5",
        x"B8",
        x"85",
        x"FF",
        x"A9",
        x"6F",
        x"03",
        x"20",
        x"72",
        x"16",
        x"4C",
        x"00",
        x"A9",
        x"25",
        x"85",
        x"20",
        x"A0",
        x"E0",
        x"A9",
        x"2B",
        x"85",
        x"2A",
        x"84",
        x"0A",
        x"A9",
        x"7F",
        x"A0",
        x"20",
        x"A2",
        x"73",
        x"9A",
        x"20",
        x"F3",
        x"A0",
        x"60",
        x"A2",
        x"F5",
        x"F0",
        x"CB",
        x"A5",
        x"73",
        x"9A",
        x"4C",
        x"E7",
        x"A0",
        x"60",
        x"A2",
        x"B5",
        x"D0",
        x"DF",
        x"A0",
        x"C1",
        x"D0",
        x"0A",
        x"A9",
        x"00",
        x"A0",
        x"06",
        x"10",
        x"B5",
        x"A5",
        x"6E",
        x"D3",
        x"20",
        x"73",
        x"D5",
        x"20",
        x"03",
        x"D0",
        x"73",
        x"E8",
        x"20",
        x"7B",
        x"A4",
        x"4C",
        x"0A",
        x"A2",
        x"AA",
        x"86",
        x"A3",
        x"A6",
        x"2C",
        x"E3",
        x"A6",
        x"03",
        x"D0",
        x"B8",
        x"A5",
        x"73",
        x"9A",
        x"20",
        x"D1",
        x"D0",
        x"61",
        x"A2",
        x"76",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"69",
        x"A0",
        x"61",
        x"A2",
        x"59",
        x"F0",
        x"00",
        x"A0",
        x"20",
        x"A9",
        x"2B",
        x"85",
        x"2A",
        x"84",
        x"0A",
        x"A9",
        x"51",
        x"A0",
        x"5F",
        x"D0",
        x"09",
        x"A9",
        x"8E",
        x"A0",
        x"06",
        x"30",
        x"B5",
        x"A5",
        x"6E",
        x"D0",
        x"20",
        x"61",
        x"A0",
        x"61",
        x"A2",
        x"73",
        x"9A",
        x"4C",
        x"57",
        x"A0",
        x"61",
        x"A2",
        x"73",
        x"9A",
        x"20",
        x"3C",
        x"A0",
        x"61",
        x"A2",
        x"07",
        x"F0",
        x"B5",
        x"A5",
        x"73",
        x"9A",
        x"20",
        x"4A",
        x"A0",
        x"61",
        x"A2",
        x"1D",
        x"D0",
        x"61",
        x"A2",
        x"42",
        x"A0",
        x"1C",
        x"D0",
        x"61",
        x"A2",
        x"2B",
        x"A0",
        x"6F",
        x"14",
        x"20",
        x"2C",
        x"A2",
        x"09",
        x"A9",
        x"72",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"10",
        x"A0",
        x"61",
        x"A2",
        x"10",
        x"30",
        x"CC",
        x"A6",
        x"73",
        x"9A",
        x"20",
        x"FC",
        x"A0",
        x"60",
        x"A2",
        x"60",
        x"00",
        x"A9",
        x"09",
        x"B5",
        x"8D",
        x"AA",
        x"A9",
        x"D4",
        x"D0",
        x"0A",
        x"C0",
        x"C8",
        x"C8",
        x"2F",
        x"A4",
        x"70",
        x"A3",
        x"20",
        x"09",
        x"95",
        x"8D",
        x"09",
        x"B5",
        x"8D",
        x"09",
        x"D5",
        x"8D",
        x"70",
        x"94",
        x"20",
        x"09",
        x"95",
        x"8D",
        x"A0",
        x"A9",
        x"6F",
        x"14",
        x"20",
        x"0B",
        x"A2",
        x"09",
        x"A9",
        x"B5",
        x"A0",
        x"AB",
        x"85",
        x"6C",
        x"25",
        x"B9",
        x"2F",
        x"84",
        x"00",
        x"A0",
        x"6F",
        x"03",
        x"20",
        x"EE",
        x"10",
        x"CA",
        x"CA",
        x"5D",
        x"A6",
        x"73",
        x"9A",
        x"20",
        x"AA",
        x"6E",
        x"06",
        x"BD",
        x"6E",
        x"05",
        x"BC",
        x"5D",
        x"86",
        x"0C",
        x"A2",
        x"E0",
        x"D0",
        x"C0",
        x"A5",
        x"61",
        x"CF",
        x"61",
        x"CA",
        x"61",
        x"B6",
        x"61",
        x"B1",
        x"61",
        x"A0",
        x"61",
        x"8A",
        x"61",
        x"80",
        x"F7",
        x"D0",
        x"CE",
        x"A0",
        x"60",
        x"A2",
        x"73",
        x"9A",
        x"4C",
        x"97",
        x"A0",
        x"60",
        x"A2",
        x"60",
        x"01",
        x"D0",
        x"C9",
        x"A5",
        x"73",
        x"9A",
        x"20",
        x"B5",
        x"A0",
        x"60",
        x"A2",
        x"E4",
        x"D0",
        x"28",
        x"91",
        x"C8",
        x"28",
        x"91",
        x"20",
        x"A0",
        x"28",
        x"91",
        x"C8",
        x"28",
        x"91",
        x"A8",
        x"00",
        x"A9",
        x"60",
        x"EE",
        x"D0",
        x"24",
        x"C6",
        x"74",
        x"7A",
        x"20",
        x"74",
        x"7A",
        x"20",
        x"74",
        x"16",
        x"20",
        x"25",
        x"A5",
        x"10",
        x"30",
        x"CA",
        x"23",
        x"A6",
        x"25",
        x"85",
        x"24",
        x"86",
        x"05",
        x"A2",
        x"29",
        x"86",
        x"28",
        x"84",
        x"4C",
        x"A9",
        x"0B",
        x"A2",
        x"7E",
        x"A0",
        x"23",
        x"86",
        x"CA",
        x"A4",
        x"A6",
        x"0B",
        x"D0",
        x"48",
        x"A9",
        x"09",
        x"A2",
        x"60",
        x"A0",
        x"23",
        x"85",
        x"A4",
        x"E5",
        x"38",
        x"86",
        x"A9",
        x"0F",
        x"10",
        x"B5",
        x"24",
        x"A4",
        x"E6",
        x"5C",
        x"85",
        x"49",
        x"A9",
        x"9F",
        x"85",
        x"80",
        x"A9",
        x"60",
        x"28",
        x"91",
        x"CF",
        x"A9",
        x"FA",
        x"D0",
        x"CA",
        x"74",
        x"7A",
        x"20",
        x"06",
        x"F0",
        x"AA",
        x"C8",
        x"01",
        x"90",
        x"00",
        x"A0",
        x"4A",
        x"01",
        x"E9",
        x"38",
        x"6D",
        x"27",
        x"20",
        x"F7",
        x"30",
        x"B5",
        x"24",
        x"0A",
        x"10",
        x"6D",
        x"32",
        x"20",
        x"60",
        x"E8",
        x"D0",
        x"CA",
        x"74",
        x"7A",
        x"20",
        x"F0",
        x"90",
        x"02",
        x"C0",
        x"C8",
        x"28",
        x"91",
        x"24",
        x"A5",
        x"2C",
        x"25",
        x"A5",
        x"03",
        x"30",
        x"26",
        x"C6",
        x"00",
        x"A0",
        x"0A",
        x"A2",
        x"25",
        x"86",
        x"24",
        x"84",
        x"26",
        x"85",
        x"CE",
        x"A0",
        x"CF",
        x"A2",
        x"6D",
        x"27",
        x"20",
        x"07",
        x"D0",
        x"FF",
        x"A0",
        x"FE",
        x"A2",
        x"6D",
        x"32",
        x"20",
        x"60",
        x"A7",
        x"E5",
        x"38",
        x"14",
        x"A9",
        x"28",
        x"84",
        x"29",
        x"86",
        x"80",
        x"A0",
        x"0B",
        x"A2",
        x"60",
        x"A7",
        x"A5",
        x"28",
        x"84",
        x"29",
        x"86",
        x"9E",
        x"A0",
        x"09",
        x"A2",
        x"60",
        x"FC",
        x"D0",
        x"8A",
        x"A5",
        x"73",
        x"9A",
        x"20",
        x"6C",
        x"2E",
        x"20",
        x"74",
        x"05",
        x"20",
        x"2E",
        x"85",
        x"00",
        x"A9",
        x"07",
        x"70",
        x"13",
        x"24",
        x"8A",
        x"85",
        x"06",
        x"A9",
        x"60",
        x"28",
        x"91",
        x"00",
        x"A9",
        x"04",
        x"90",
        x"60",
        x"C9",
        x"04",
        x"90",
        x"11",
        x"C9",
        x"28",
        x"B1",
        x"72",
        x"BE",
        x"4C",
        x"6F",
        x"EF",
        x"20",
        x"6E",
        x"E3",
        x"20",
        x"6D",
        x"40",
        x"20",
        x"6D",
        x"A2",
        x"20",
        x"70",
        x"EA",
        x"20",
        x"6C",
        x"4E",
        x"20",
        x"70",
        x"97",
        x"20",
        x"90",
        x"85",
        x"80",
        x"A9",
        x"73",
        x"58",
        x"20",
        x"6E",
        x"A4",
        x"20",
        x"0A",
        x"30",
        x"90",
        x"24",
        x"6E",
        x"C3",
        x"20",
        x"6C",
        x"4E",
        x"20",
        x"6F",
        x"DF",
        x"20",
        x"6F",
        x"B5",
        x"20",
        x"AF",
        x"10",
        x"B5",
        x"24",
        x"72",
        x"8E",
        x"20",
        x"6F",
        x"C9",
        x"20",
        x"72",
        x"BE",
        x"4C",
        x"72",
        x"B8",
        x"4C",
        x"03",
        x"D0",
        x"B5",
        x"A5",
        x"6F",
        x"E9",
        x"20",
        x"6E",
        x"E8",
        x"20",
        x"6D",
        x"49",
        x"20",
        x"6D",
        x"B1",
        x"20",
        x"70",
        x"EA",
        x"20",
        x"6C",
        x"45",
        x"20",
        x"70",
        x"97",
        x"20",
        x"90",
        x"85",
        x"80",
        x"A9",
        x"73",
        x"0E",
        x"20",
        x"6E",
        x"85",
        x"20",
        x"0A",
        x"30",
        x"90",
        x"24",
        x"6E",
        x"8B",
        x"20",
        x"6C",
        x"45",
        x"20",
        x"0D",
        x"F0",
        x"B8",
        x"A5",
        x"6F",
        x"DF",
        x"20",
        x"6C",
        x"8B",
        x"4C",
        x"6F",
        x"DC",
        x"20",
        x"06",
        x"D0",
        x"B5",
        x"A5",
        x"6F",
        x"B5",
        x"20",
        x"6F",
        x"CC",
        x"20",
        x"72",
        x"94",
        x"20",
        x"4D",
        x"D0",
        x"B5",
        x"A5",
        x"70",
        x"9A",
        x"20",
        x"0D",
        x"F0",
        x"72",
        x"8E",
        x"20",
        x"6F",
        x"C9",
        x"20",
        x"62",
        x"F0",
        x"72",
        x"94",
        x"20",
        x"6F",
        x"CC",
        x"20",
        x"08",
        x"F0",
        x"B5",
        x"A5",
        x"70",
        x"9A",
        x"20",
        x"71",
        x"B6",
        x"4C",
        x"6D",
        x"FF",
        x"20",
        x"70",
        x"06",
        x"20",
        x"71",
        x"96",
        x"4C",
        x"6D",
        x"EC",
        x"20",
        x"70",
        x"06",
        x"20",
        x"60",
        x"60",
        x"A2",
        x"AF",
        x"A0",
        x"04",
        x"D0",
        x"60",
        x"A2",
        x"A9",
        x"A0",
        x"06",
        x"30",
        x"0C",
        x"D0",
        x"60",
        x"A2",
        x"A3",
        x"A0",
        x"06",
        x"D0",
        x"B5",
        x"A5",
        x"80",
        x"00",
        x"30",
        x"00",
        x"15",
        x"00",
        x"06",
        x"00",
        x"03",
        x"68",
        x"6C",
        x"4C",
        x"0C",
        x"0F",
        x"8D",
        x"00",
        x"A9",
        x"E1",
        x"F0",
        x"C0",
        x"A5",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"E0",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"D9",
        x"A0",
        x"F3",
        x"D0",
        x"B8",
        x"A5",
        x"68",
        x"AF",
        x"4C",
        x"73",
        x"9A",
        x"20",
        x"6C",
        x"2E",
        x"20",
        x"03",
        x"D0",
        x"60",
        x"A2",
        x"9D",
        x"A0",
        x"09",
        x"D0",
        x"60",
        x"A2",
        x"97",
        x"A0",
        x"06",
        x"30",
        x"11",
        x"D0",
        x"60",
        x"A2",
        x"91",
        x"A0",
        x"06",
        x"D0",
        x"B5",
        x"A5",
        x"18",
        x"F0",
        x"10",
        x"29",
        x"8B",
        x"A5",
        x"2B",
        x"F0",
        x"B8",
        x"A5",
        x"7D",
        x"43",
        x"4C",
        x"03",
        x"30",
        x"0C",
        x"0F",
        x"2C",
        x"74",
        x"05",
        x"20",
        x"2E",
        x"84",
        x"00",
        x"A0",
        x"02",
        x"F0",
        x"20",
        x"29",
        x"8B",
        x"A5",
        x"04",
        x"A0",
        x"42",
        x"D0",
        x"13",
        x"A5",
        x"57",
        x"66",
        x"02",
        x"90",
        x"9A",
        x"C5",
        x"8E",
        x"A5",
        x"08",
        x"B0",
        x"99",
        x"C5",
        x"A5",
        x"A5",
        x"0E",
        x"B0",
        x"14",
        x"C9",
        x"A6",
        x"A5",
        x"71",
        x"53",
        x"20",
        x"26",
        x"84",
        x"C8",
        x"C8",
        x"07",
        x"D0",
        x"3C",
        x"C9",
        x"05",
        x"F0",
        x"28",
        x"C9",
        x"0A",
        x"F0",
        x"14",
        x"C9",
        x"91",
        x"A5",
        x"01",
        x"A0",
        x"17",
        x"D0",
        x"92",
        x"A5",
        x"92",
        x"E6",
        x"02",
        x"D0",
        x"91",
        x"E6",
        x"8F",
        x"E6",
        x"8E",
        x"E6",
        x"8D",
        x"85",
        x"00",
        x"A9",
        x"0E",
        x"90",
        x"3C",
        x"C9",
        x"8D",
        x"A5",
        x"68",
        x"A1",
        x"4C",
        x"6C",
        x"57",
        x"20",
        x"90",
        x"85",
        x"00",
        x"A9",
        x"71",
        x"22",
        x"20",
        x"0C",
        x"0F",
        x"8D",
        x"00",
        x"A9",
        x"6D",
        x"0D",
        x"20",
        x"15",
        x"90",
        x"14",
        x"C9",
        x"A7",
        x"A5",
        x"6A",
        x"47",
        x"4C",
        x"03",
        x"F0",
        x"13",
        x"A5",
        x"22",
        x"D0",
        x"14",
        x"A5",
        x"71",
        x"D4",
        x"20",
        x"03",
        x"D0",
        x"71",
        x"DC",
        x"20",
        x"08",
        x"D0",
        x"71",
        x"EC",
        x"20",
        x"0A",
        x"10",
        x"07",
        x"F0",
        x"B5",
        x"A5",
        x"02",
        x"A2",
        x"71",
        x"E2",
        x"20",
        x"03",
        x"D0",
        x"71",
        x"FA",
        x"20",
        x"05",
        x"10",
        x"B5",
        x"24",
        x"F9",
        x"10",
        x"CA",
        x"C3",
        x"95",
        x"A0",
        x"B5",
        x"F5",
        x"F0",
        x"15",
        x"90",
        x"C3",
        x"D5",
        x"A0",
        x"B5",
        x"1B",
        x"30",
        x"CA",
        x"03",
        x"A2",
        x"6D",
        x"94",
        x"20",
        x"03",
        x"90",
        x"CC",
        x"C5",
        x"A1",
        x"A5",
        x"09",
        x"30",
        x"9F",
        x"A5",
        x"54",
        x"85",
        x"53",
        x"85",
        x"00",
        x"A9",
        x"D8",
        x"F7",
        x"D0",
        x"E8",
        x"A3",
        x"95",
        x"A3",
        x"75",
        x"56",
        x"B5",
        x"FD",
        x"A2",
        x"18",
        x"F8",
        x"56",
        x"F0",
        x"54",
        x"05",
        x"53",
        x"A5",
        x"68",
        x"A1",
        x"4C",
        x"6C",
        x"6E",
        x"20",
        x"B5",
        x"86",
        x"FF",
        x"A2",
        x"02",
        x"10",
        x"CD",
        x"24",
        x"7F",
        x"A2",
        x"08",
        x"D0",
        x"B5",
        x"A5",
        x"00",
        x"A2",
        x"B4",
        x"85",
        x"68",
        x"6C",
        x"4C",
        x"70",
        x"9A",
        x"20",
        x"6F",
        x"CC",
        x"20",
        x"03",
        x"30",
        x"6F",
        x"C9",
        x"20",
        x"05",
        x"D0",
        x"B5",
        x"A5",
        x"12",
        x"D0",
        x"C0",
        x"C9",
        x"B4",
        x"05",
        x"4A",
        x"01",
        x"F0",
        x"B5",
        x"A4",
        x"80",
        x"A9",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"E0",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"D9",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"3C",
        x"A0",
        x"07",
        x"F0",
        x"B5",
        x"A4",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"4A",
        x"A0",
        x"1D",
        x"D0",
        x"61",
        x"A2",
        x"EE",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"E7",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"69",
        x"A0",
        x"14",
        x"10",
        x"B5",
        x"24",
        x"68",
        x"A1",
        x"4C",
        x"6C",
        x"57",
        x"20",
        x"5F",
        x"F0",
        x"B4",
        x"A5",
        x"A5",
        x"85",
        x"00",
        x"A9",
        x"90",
        x"85",
        x"00",
        x"A9",
        x"71",
        x"22",
        x"20",
        x"07",
        x"90",
        x"14",
        x"C9",
        x"A6",
        x"85",
        x"A7",
        x"A5",
        x"1D",
        x"F0",
        x"A4",
        x"C6",
        x"21",
        x"70",
        x"13",
        x"24",
        x"76",
        x"F0",
        x"B8",
        x"A5",
        x"70",
        x"94",
        x"20",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"E0",
        x"A0",
        x"73",
        x"9A",
        x"20",
        x"61",
        x"A2",
        x"D9",
        x"A0",
        x"0E",
        x"D0",
        x"B8",
        x"A5",
        x"0C",
        x"0F",
        x"8D",
        x"00",
        x"A9",
        x"6D",
        x"0D",
        x"20",
        x"69",
        x"1B",
        x"4C",
        x"8E",
        x"86",
        x"6D",
        x"76",
        x"20",
        x"A7",
        x"E6",
        x"A5",
        x"C6",
        x"76",
        x"34",
        x"20",
        x"6C",
        x"25",
        x"BD",
        x"03",
        x"D0",
        x"80",
        x"A9",
        x"76",
        x"34",
        x"20",
        x"80",
        x"A9",
        x"09",
        x"D0",
        x"0A",
        x"E0",
        x"28",
        x"91",
        x"01",
        x"69",
        x"18",
        x"20",
        x"A0",
        x"28",
        x"91",
        x"00",
        x"A0",
        x"60",
        x"09",
        x"2C",
        x"70",
        x"09",
        x"03",
        x"10",
        x"B5",
        x"24",
        x"AA",
        x"48",
        x"B5",
        x"73",
        x"C6",
        x"20",
        x"3B",
        x"95",
        x"3C",
        x"F6",
        x"02",
        x"90",
        x"21",
        x"69",
        x"3B",
        x"B5",
        x"18",
        x"69",
        x"5B",
        x"4C",
        x"74",
        x"05",
        x"20",
        x"2E",
        x"85",
        x"EC",
        x"A9",
        x"07",
        x"F0",
        x"40",
        x"29",
        x"0E",
        x"10",
        x"48",
        x"B5",
        x"24",
        x"A6",
        x"EE",
        x"D0",
        x"23",
        x"C6",
        x"74",
        x"6E",
        x"20",
        x"F7",
        x"10",
        x"88",
        x"E8",
        x"28",
        x"91",
        x"02",
        x"00",
        x"BD",
        x"03",
        x"A0",
        x"74",
        x"64",
        x"20",
        x"69",
        x"1D",
        x"4C",
        x"DF",
        x"F0",
        x"60",
        x"C9",
        x"07",
        x"F0",
        x"24",
        x"C9",
        x"CA",
        x"F0",
        x"1B",
        x"C9",
        x"D1",
        x"F0",
        x"12",
        x"C9",
        x"D2",
        x"F0",
        x"09",
        x"C9",
        x"69",
        x"59",
        x"4C",
        x"6C",
        x"FE",
        x"20",
        x"20",
        x"A0",
        x"6C",
        x"FE",
        x"20",
        x"00",
        x"A0",
        x"69",
        x"1B",
        x"4C",
        x"EF",
        x"D0",
        x"23",
        x"C6",
        x"74",
        x"6E",
        x"20",
        x"F8",
        x"10",
        x"88",
        x"E8",
        x"AA",
        x"28",
        x"91",
        x"8A",
        x"03",
        x"A0",
        x"23",
        x"84",
        x"04",
        x"A0",
        x"30",
        x"A2",
        x"2C",
        x"20",
        x"A2",
        x"69",
        x"18",
        x"4C",
        x"18",
        x"A9",
        x"28",
        x"85",
        x"29",
        x"C6",
        x"02",
        x"B0",
        x"5F",
        x"E9",
        x"28",
        x"A5",
        x"38",
        x"ED",
        x"D0",
        x"23",
        x"C6",
        x"74",
        x"6E",
        x"20",
        x"F6",
        x"10",
        x"88",
        x"E8",
        x"02",
        x"00",
        x"9D",
        x"74",
        x"2C",
        x"20",
        x"03",
        x"A0",
        x"74",
        x"64",
        x"20",
        x"73",
        x"C6",
        x"20",
        x"3B",
        x"95",
        x"3C",
        x"D6",
        x"02",
        x"B0",
        x"21",
        x"E9",
        x"3B",
        x"B5",
        x"38",
        x"5E",
        x"D0",
        x"BC",
        x"F0",
        x"47",
        x"94",
        x"3C",
        x"94",
        x"00",
        x"A0",
        x"24",
        x"A6",
        x"28",
        x"91",
        x"02",
        x"60",
        x"BD",
        x"C8",
        x"E8",
        x"28",
        x"91",
        x"02",
        x"60",
        x"BD",
        x"E8",
        x"20",
        x"A0",
        x"28",
        x"91",
        x"02",
        x"60",
        x"BD",
        x"C8",
        x"E8",
        x"28",
        x"91",
        x"02",
        x"60",
        x"BD",
        x"00",
        x"A0",
        x"AA",
        x"0A",
        x"8A",
        x"E4",
        x"D0",
        x"1B",
        x"C9",
        x"F4",
        x"F0",
        x"12",
        x"C9",
        x"F5",
        x"F0",
        x"09",
        x"C9",
        x"EB",
        x"D0",
        x"1C",
        x"A9",
        x"AC",
        x"18",
        x"A9",
        x"6A",
        x"FC",
        x"4C",
        x"C1",
        x"10",
        x"CA",
        x"CA",
        x"47",
        x"F6",
        x"24",
        x"A6",
        x"74",
        x"16",
        x"20",
        x"14",
        x"A9",
        x"02",
        x"60",
        x"9D",
        x"74",
        x"55",
        x"20",
        x"02",
        x"60",
        x"9D",
        x"74",
        x"56",
        x"20",
        x"20",
        x"A0",
        x"02",
        x"60",
        x"9D",
        x"74",
        x"55",
        x"20",
        x"02",
        x"60",
        x"9D",
        x"74",
        x"57",
        x"20",
        x"00",
        x"A0",
        x"AA",
        x"0A",
        x"8A",
        x"36",
        x"D0",
        x"7F",
        x"29",
        x"70",
        x"10",
        x"24",
        x"86",
        x"47",
        x"B5",
        x"73",
        x"C4",
        x"20",
        x"14",
        x"E6",
        x"37",
        x"F0",
        x"3C",
        x"B5",
        x"0A",
        x"A2",
        x"14",
        x"85",
        x"00",
        x"A9",
        x"0C",
        x"09",
        x"8E",
        x"00",
        x"A2",
        x"02",
        x"D0",
        x"08",
        x"29",
        x"01",
        x"A2",
        x"5C",
        x"A5",
        x"5C",
        x"C6",
        x"0F",
        x"F0",
        x"5C",
        x"A5",
        x"0C",
        x"0C",
        x"8E",
        x"03",
        x"D0",
        x"5A",
        x"A5",
        x"0C",
        x"0D",
        x"8E",
        x"03",
        x"D0",
        x"59",
        x"A5",
        x"00",
        x"A2",
        x"5A",
        x"C6",
        x"59",
        x"C6",
        x"2C",
        x"85",
        x"FA",
        x"F0",
        x"2C",
        x"C5",
        x"8B",
        x"A5",
        x"5E",
        x"86",
        x"FF",
        x"A2",
        x"0C",
        x"0F",
        x"8E",
        x"01",
        x"A2",
        x"0C",
        x"0A",
        x"8E",
        x"00",
        x"A2",
        x"2C",
        x"01",
        x"A2",
        x"71",
        x"2A",
        x"20",
        x"06",
        x"D0",
        x"B8",
        x"A5",
        x"6C",
        x"78",
        x"20",
        x"6F",
        x"C9",
        x"20",
        x"73",
        x"54",
        x"20",
        x"71",
        x"27",
        x"20",
        x"6F",
        x"23",
        x"20",
        x"6E",
        x"64",
        x"20",
        x"6C",
        x"45",
        x"20",
        x"09",
        x"F0",
        x"6E",
        x"13",
        x"20",
        x"6C",
        x"45",
        x"20",
        x"08",
        x"F0",
        x"CB",
        x"A5",
        x"58",
        x"A4",
        x"85",
        x"CA",
        x"A5",
        x"C7",
        x"E6",
        x"6F",
        x"B2",
        x"20",
        x"68",
        x"00",
        x"20",
        x"6F",
        x"96",
        x"20",
        x"60",
        x"F5",
        x"10",
        x"0C",
        x"0F",
        x"2C",
        x"70",
        x"85",
        x"20",
        x"70",
        x"26",
        x"20",
        x"6F",
        x"B2",
        x"20",
        x"6F",
        x"96",
        x"20",
        x"AC",
        x"F0",
        x"70",
        x"82",
        x"20",
        x"7E",
        x"A1",
        x"20",
        x"0C",
        x"08",
        x"99",
        x"00",
        x"A9",
        x"2C",
        x"01",
        x"A9",
        x"A8",
        x"01",
        x"29",
        x"98",
        x"07",
        x"30",
        x"0C",
        x"07",
        x"2C",
        x"00",
        x"A0",
        x"F3",
        x"10",
        x"88",
        x"0A",
        x"10",
        x"0C",
        x"05",
        x"B9",
        x"0F",
        x"10",
        x"0C",
        x"0D",
        x"B9",
        x"01",
        x"A0",
        x"E1",
        x"D0",
        x"B5",
        x"C6",
        x"04",
        x"30",
        x"B5",
        x"A5",
        x"1E",
        x"F0",
        x"77",
        x"75",
        x"20",
        x"01",
        x"A0",
        x"25",
        x"90",
        x"7C",
        x"F8",
        x"20",
        x"79",
        x"A2",
        x"20",
        x"0C",
        x"01",
        x"8D",
        x"0C",
        x"00",
        x"8D",
        x"01",
        x"A9",
        x"49",
        x"30",
        x"0C",
        x"0F",
        x"2C",
        x"7B",
        x"B8",
        x"20",
        x"6F",
        x"A1",
        x"20",
        x"58",
        x"54",
        x"09",
        x"58",
        x"30",
        x"31",
        x"53",
        x"4D",
        x"0D",
        x"3B",
        x"0D",
        x"53",
        x"54",
        x"52",
        x"09",
        x"32",
        x"30",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"0D",
        x"30",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"41",
        x"44",
        x"4C",
        x"09",
        x"0D",
        x"32",
        x"30",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"53",
        x"43",
        x"42",
        x"09",
        x"0D",
        x"48",
        x"30",
        x"39",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"50",
        x"4D",
        x"43",
        x"09",
        x"0D",
        x"32",
        x"30",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"43",
        x"43",
        x"42",
        x"09",
        x"0D",
        x"48",
        x"31",
        x"31",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"50",
        x"4D",
        x"43",
        x"09",
        x"0D",
        x"4C",
        x"44",
        x"41",
        x"46",
        x"55",
        x"42",
        x"4D",
        x"3A",
        x"59",
        x"49",
        x"09",
        x"41",
        x"44",
        x"4C",
        x"09",
        x"31",
        x"4E",
        x"45",
        x"54",
        x"53",
        x"4D",
        x"0D",
        x"58",
        x"4E",
        x"49",
        x"09",
        x"34",
        x"30",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"0D",
        x"59",
        x"4E",
        x"49",
        x"09",
        x"33",
        x"30",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"0D",
        x"53",
        x"54",
        x"52",
        x"09",
        x"0D",
        x"48",
        x"30",
        x"31",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"41",
        x"44",
        x"4C",
        x"09",
        x"38",
        x"32",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"0D",
        x"31",
        x"4E",
        x"45",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"45",
        x"4E",
        x"42",
        x"09",
        x"0D",
        x"48",
        x"44",
        x"31",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"50",
        x"4D",
        x"43",
        x"09",
        x"0D",
        x"38",
        x"32",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"51",
        x"45",
        x"42",
        x"09",
        x"0D",
        x"32",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"50",
        x"4D",
        x"43",
        x"09",
        x"0D",
        x"48",
        x"46",
        x"31",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"44",
        x"4E",
        x"41",
        x"09",
        x"0D",
        x"4C",
        x"44",
        x"41",
        x"46",
        x"55",
        x"42",
        x"4D",
        x"3A",
        x"20",
        x"5A",
        x"09",
        x"43",
        x"44",
        x"41",
        x"09",
        x"0D",
        x"43",
        x"4C",
        x"43",
        x"09",
        x"0D",
        x"41",
        x"59",
        x"54",
        x"09",
        x"31",
        x"32",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"0D",
        x"38",
        x"32",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"43",
        x"43",
        x"42",
        x"09",
        x"0D",
        x"48",
        x"45",
        x"35",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"50",
        x"4D",
        x"43",
        x"09",
        x"0D",
        x"4C",
        x"44",
        x"41",
        x"46",
        x"55",
        x"42",
        x"4D",
        x"3A",
        x"20",
        x"5A",
        x"09",
        x"41",
        x"44",
        x"4C",
        x"09",
        x"0D",
        x"31",
        x"32",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"45",
        x"4E",
        x"42",
        x"09",
        x"0D",
        x"38",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"50",
        x"4D",
        x"43",
        x"09",
        x"32",
        x"31",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"0D",
        x"38",
        x"32",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"53",
        x"43",
        x"42",
        x"09",
        x"0D",
        x"31",
        x"32",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"43",
        x"43",
        x"42",
        x"09",
        x"0D",
        x"48",
        x"32",
        x"41",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"50",
        x"4D",
        x"43",
        x"09",
        x"0D",
        x"4C",
        x"44",
        x"41",
        x"46",
        x"55",
        x"42",
        x"4D",
        x"3A",
        x"20",
        x"5A",
        x"09",
        x"41",
        x"44",
        x"4C",
        x"09",
        x"0D",
        x"32",
        x"31",
        x"31",
        x"54",
        x"53",
        x"4D",
        x"3A",
        x"20",
        x"52",
        x"09",
        x"45",
        x"4E",
        x"42",
        x"09",
        x"0D",
        x"48",
        x"42",
        x"2F",
        x"20",
        x"49",
        x"09",
        x"50",
        x"4D",
        x"43",
        x"09",
        x"0D",
        x"48",
        x"44",
        x"41",
        x"46",
        x"55",
        x"42",
        x"4D",
        x"3A",
        x"20",
        x"5A",
        x"09",
        x"41",
        x"44",
        x"4C",
        x"09",
        x"30",
        x"4E",
        x"45",
        x"54",
        x"53",
        x"4D",
        x"0D",
        x"3B",
        x"0D",
        x"53",
        x"54",
        x"52",
        x"09",
        x"0D",
        x"4C",
        x"44",
        x"41",
        x"46",
        x"55",
        x"42",
        x"4D",
        x"3A",
        x"59",
        x"49",
        x"09",
        x"09",
        x"86",
        x"02",
        x"09",
        x"E3",
        x"03",
        x"01",
        x"03",
        x"00",
        x"08",
        x"9B",
        x"0B",
        x"7B",
        x"B5",
        x"A9",
        x"0A",
        x"58",
        x"03",
        x"09",
        x"FB",
        x"02",
        x"00",
        x"02",
        x"01",
        x"0B",
        x"64",
        x"08",
        x"84",
        x"B5",
        x"A9",
        x"09",
        x"08",
        x"03",
        x"80",
        x"07",
        x"06",
        x"02",
        x"80",
        x"09",
        x"07",
        x"04",
        x"80",
        x"08",
        x"06",
        x"05",
        x"80",
        x"00",
        x"08",
        x"00",
        x"06",
        x"05",
        x"00",
        x"08",
        x"06",
        x"05",
        x"09",
        x"00",
        x"07",
        x"00",
        x"00",
        x"04",
        x"09",
        x"07",
        x"04",
        x"09",
        x"08",
        x"00",
        x"00",
        x"08",
        x"09",
        x"03",
        x"00",
        x"03",
        x"00",
        x"00",
        x"07",
        x"06",
        x"06",
        x"07",
        x"00",
        x"02",
        x"02",
        x"01",
        x"00",
        x"01",
        x"00",
        x"00",
        x"01",
        x"01",
        x"01",
        x"01",
        x"00",
        x"01",
        x"00",
        x"01",
        x"01",
        x"00",
        x"01",
        x"01",
        x"01",
        x"00",
        x"00",
        x"01",
        x"01",
        x"01",
        x"01",
        x"00",
        x"01",
        x"01",
        x"01",
        x"01",
        x"00",
        x"00",
        x"01",
        x"01",
        x"01",
        x"00",
        x"01",
        x"C8",
        x"F0",
        x"C8",
        x"F0",
        x"E0",
        x"E8",
        x"F0",
        x"F4",
        x"F0",
        x"F0",
        x"F0",
        x"F0",
        x"02",
        x"02",
        x"02",
        x"02",
        x"04",
        x"03",
        x"02",
        x"01",
        x"03",
        x"01",
        x"03",
        x"01",
        x"01",
        x"02",
        x"02",
        x"03",
        x"F4",
        x"C8",
        x"A8",
        x"80",
        x"B0",
        x"90",
        x"70",
        x"60",
        x"90",
        x"70",
        x"60",
        x"40",
        x"60",
        x"40",
        x"40",
        x"20",
        x"A0",
        x"80",
        x"80",
        x"50",
        x"A0",
        x"60",
        x"80",
        x"40",
        x"50",
        x"30",
        x"30",
        x"50",
        x"60",
        x"30",
        x"20",
        x"20",
        x"01",
        x"02",
        x"01",
        x"02",
        x"01",
        x"01",
        x"01",
        x"01",
        x"01",
        x"01",
        x"02",
        x"02",
        x"01",
        x"02",
        x"02",
        x"03",
        x"07",
        x"07",
        x"07",
        x"07",
        x"07",
        x"07",
        x"06",
        x"05",
        x"06",
        x"06",
        x"05",
        x"04",
        x"05",
        x"05",
        x"04",
        x"03",
        x"00",
        x"00",
        x"03",
        x"02",
        x"02",
        x"03",
        x"02",
        x"01",
        x"00",
        x"00",
        x"02",
        x"02",
        x"03",
        x"03",
        x"02",
        x"02",
        x"00",
        x"00",
        x"02",
        x"02",
        x"02",
        x"02",
        x"02",
        x"01",
        x"00",
        x"00",
        x"02",
        x"02",
        x"02",
        x"02",
        x"02",
        x"01",
        x"00",
        x"00",
        x"02",
        x"02",
        x"03",
        x"03",
        x"02",
        x"02",
        x"00",
        x"00",
        x"02",
        x"02",
        x"02",
        x"02",
        x"02",
        x"00",
        x"00",
        x"00",
        x"02",
        x"02",
        x"02",
        x"02",
        x"02",
        x"00",
        x"00",
        x"00",
        x"01",
        x"03",
        x"01",
        x"02",
        x"01",
        x"02",
        x"00",
        x"00",
        x"01",
        x"03",
        x"02",
        x"01",
        x"01",
        x"00",
        x"00",
        x"00",
        x"01",
        x"03",
        x"02",
        x"01",
        x"01",
        x"00",
        x"00",
        x"00",
        x"03",
        x"02",
        x"02",
        x"03",
        x"02",
        x"02",
        x"00",
        x"00",
        x"02",
        x"02",
        x"03",
        x"03",
        x"02",
        x"02",
        x"00",
        x"00",
        x"02",
        x"02",
        x"02",
        x"02",
        x"02",
        x"01",
        x"00",
        x"00",
        x"02",
        x"02",
        x"02",
        x"02",
        x"02",
        x"01",
        x"00",
        x"00",
        x"01",
        x"03",
        x"01",
        x"02",
        x"01",
        x"02",
        x"00",
        x"00",
        x"01",
        x"03",
        x"02",
        x"01",
        x"01",
        x"00",
        x"00",
        x"00",
        x"01",
        x"03",
        x"02",
        x"01",
        x"01",
        x"00",
        x"00",
        x"00",
        x"00",
        x"03",
        x"00",
        x"02",
        x"03",
        x"02",
        x"00",
        x"00",
        x"00",
        x"01",
        x"01",
        x"00",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"3C",
        x"CF",
        x"CC",
        x"F0",
        x"3C",
        x"33",
        x"03",
        x"00",
        x"0C",
        x"00",
        x"00",
        x"30",
        x"00",
        x"FC",
        x"CC",
        x"FF",
        x"F0",
        x"33",
        x"FF",
        x"03",
        x"C0",
        x"00",
        x"00",
        x"00",
        x"03",
        x"00",
        x"FC",
        x"FC",
        x"1F",
        x"F0",
        x"F3",
        x"7F",
        x"0E",
        x"00",
        x"00",
        x"08",
        x"00",
        x"00",
        x"20",
        x"FC",
        x"F3",
        x"9F",
        x"F3",
        x"CF",
        x"7F",
        x"00",
        x"00",
        x"03",
        x"00",
        x"00",
        x"0C",
        x"00",
        x"CC",
        x"33",
        x"FF",
        x"30",
        x"CF",
        x"FC",
        x"C3",
        x"0C",
        x"30",
        x"00",
        x"33",
        x"C0",
        x"00",
        x"CC",
        x"3C",
        x"F3",
        x"30",
        x"F3",
        x"CC",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"3C",
        x"CF",
        x"F3",
        x"F0",
        x"3C",
        x"CF",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"3C",
        x"CF",
        x"F3",
        x"F0",
        x"3C",
        x"CF",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"3C",
        x"CF",
        x"13",
        x"F0",
        x"3C",
        x"4F",
        x"0E",
        x"00",
        x"00",
        x"09",
        x"00",
        x"00",
        x"24",
        x"3C",
        x"CF",
        x"93",
        x"F3",
        x"3C",
        x"4F",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"3C",
        x"CF",
        x"F3",
        x"F0",
        x"3C",
        x"CF",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"3C",
        x"CF",
        x"F3",
        x"F0",
        x"3C",
        x"CF",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"FE",
        x"FF",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"E0",
        x"FF",
        x"33",
        x"00",
        x"00",
        x"40",
        x"00",
        x"00",
        x"00",
        x"81",
        x"E1",
        x"3F",
        x"07",
        x"05",
        x"00",
        x"00",
        x"1C",
        x"00",
        x"00",
        x"F0",
        x"F9",
        x"7F",
        x"0E",
        x"00",
        x"02",
        x"08",
        x"00",
        x"08",
        x"20",
        x"7C",
        x"FE",
        x"9F",
        x"73",
        x"00",
        x"00",
        x"40",
        x"01",
        x"00",
        x"00",
        x"86",
        x"FF",
        x"1C",
        x"00",
        x"00",
        x"40",
        x"00",
        x"00",
        x"00",
        x"01",
        x"F8",
        x"FF",
        x"0C",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"F8",
        x"FF",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"06",
        x"00",
        x"00",
        x"18",
        x"00",
        x"FC",
        x"07",
        x"FE",
        x"F0",
        x"1F",
        x"F8",
        x"03",
        x"00",
        x"06",
        x"00",
        x"00",
        x"18",
        x"00",
        x"FC",
        x"67",
        x"FE",
        x"F0",
        x"9F",
        x"F9",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"FC",
        x"99",
        x"1F",
        x"F0",
        x"67",
        x"7E",
        x"0E",
        x"80",
        x"01",
        x"08",
        x"00",
        x"06",
        x"20",
        x"FC",
        x"99",
        x"9F",
        x"F3",
        x"67",
        x"7E",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"FC",
        x"67",
        x"FE",
        x"F0",
        x"9F",
        x"F9",
        x"03",
        x"00",
        x"06",
        x"00",
        x"00",
        x"18",
        x"00",
        x"FC",
        x"07",
        x"FE",
        x"F0",
        x"1F",
        x"F8",
        x"03",
        x"00",
        x"06",
        x"00",
        x"00",
        x"18",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"0E",
        x"00",
        x"00",
        x"08",
        x"00",
        x"00",
        x"20",
        x"00",
        x"00",
        x"80",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"9C",
        x"33",
        x"F3",
        x"70",
        x"CE",
        x"CC",
        x"C3",
        x"39",
        x"33",
        x"0F",
        x"E7",
        x"0C",
        x"00",
        x"9C",
        x"33",
        x"00",
        x"00",
        x"C0",
        x"FF",
        x"03",
        x"00",
        x"FF",
        x"0F",
        x"FF",
        x"0C",
        x"00",
        x"FC",
        x"33",
        x"00",
        x"F0",
        x"CF",
        x"4C",
        x"0E",
        x"00",
        x"30",
        x"09",
        x"00",
        x"C0",
        x"24",
        x"FC",
        x"33",
        x"93",
        x"F3",
        x"CF",
        x"00",
        x"00",
        x"00",
        x"03",
        x"00",
        x"00",
        x"CC",
        x"3C",
        x"FC",
        x"33",
        x"F3",
        x"F0",
        x"CF",
        x"CC",
        x"03",
        x"00",
        x"03",
        x"00",
        x"00",
        x"0C",
        x"00",
        x"3C",
        x"FF",
        x"FC",
        x"F0",
        x"FC",
        x"F3",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"02",
        x"00",
        x"00",
        x"08",
        x"00",
        x"3C",
        x"27",
        x"FF",
        x"F0",
        x"9C",
        x"FC",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"FC",
        x"99",
        x"FF",
        x"F0",
        x"67",
        x"FE",
        x"03",
        x"80",
        x"01",
        x"00",
        x"00",
        x"06",
        x"00",
        x"3C",
        x"FF",
        x"19",
        x"F0",
        x"FC",
        x"67",
        x"0E",
        x"80",
        x"81",
        x"09",
        x"00",
        x"06",
        x"26",
        x"FC",
        x"99",
        x"99",
        x"F3",
        x"67",
        x"06",
        x"C0",
        x"80",
        x"19",
        x"00",
        x"03",
        x"66",
        x"3E",
        x"CC",
        x"99",
        x"F9",
        x"30",
        x"67",
        x"E6",
        x"03",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"CC",
        x"27",
        x"FF",
        x"30",
        x"9F",
        x"FC",
        x"03",
        x"00",
        x"02",
        x"00",
        x"00",
        x"08",
        x"00",
        x"00",
        x"80",
        x"01",
        x"00",
        x"00",
        x"06",
        x"00",
        x"CC",
        x"99",
        x"CF",
        x"30",
        x"67",
        x"3E",
        x"C3",
        x"80",
        x"19",
        x"00",
        x"03",
        x"66",
        x"00",
        x"FC",
        x"99",
        x"F9",
        x"F0",
        x"67",
        x"E6",
        x"03",
        x"00",
        x"80",
        x"0F",
        x"00",
        x"00",
        x"00",
        x"7C",
        x"FE",
        x"01",
        x"F0",
        x"F9",
        x"67",
        x"0E",
        x"80",
        x"81",
        x"09",
        x"00",
        x"06",
        x"26",
        x"CC",
        x"99",
        x"99",
        x"33",
        x"67",
        x"06",
        x"C0",
        x"9C",
        x"19",
        x"00",
        x"70",
        x"E6",
        x"3F",
        x"C0",
        x"99",
        x"FF",
        x"30",
        x"67",
        x"00",
        x"C0",
        x"00",
        x"00",
        x"00",
        x"03",
        x"60",
        x"3E",
        x"FC",
        x"99",
        x"F9",
        x"F0",
        x"67",
        x"E6",
        x"03",
        x"80",
        x"01",
        x"00",
        x"00",
        x"06",
        x"00",
        x"62",
        x"7B",
        x"62",
        x"D0",
        x"63",
        x"25",
        x"63",
        x"7A",
        x"63",
        x"CF",
        x"64",
        x"24",
        x"64",
        x"79",
        x"64",
        x"CE",
        x"62",
        x"27",
        x"62",
        x"7C",
        x"62",
        x"D1",
        x"63",
        x"26",
        x"63",
        x"7B",
        x"63",
        x"D0",
        x"64",
        x"25",
        x"64",
        x"7A",
        x"04",
        x"00",
        x"03",
        x"04",
        x"00",
        x"01",
        x"04",
        x"05",
        x"07",
        x"04",
        x"00",
        x"01",
        x"04",
        x"03",
        x"05",
        x"04",
        x"06",
        x"07",
        x"E5",
        x"ED",
        x"E1",
        x"E7",
        x"04",
        x"09",
        x"C7",
        x"F2",
        x"E5",
        x"F6",
        x"EF",
        x"04",
        x"0A",
        x"87",
        x"BF",
        x"C6",
        x"B5",
        x"C2",
        x"04",
        x"09",
        x"D8",
        x"B7",
        x"B1",
        x"BD",
        x"B5",
        x"04",
        x"0A",
        x"98",
        x"AD",
        x"AE",
        x"AF",
        x"DC",
        x"DD",
        x"DE",
        x"DF",
        x"07",
        x"0A",
        x"59",
        x"5E",
        x"5C",
        x"02",
        x"0A",
        x"54",
        x"C4",
        x"B1",
        x"BE",
        x"BB",
        x"B0",
        x"B0",
        x"5F",
        x"5D",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"C0",
        x"C4",
        x"C3",
        x"11",
        x"0B",
        x"15",
        x"82",
        x"80",
        x"02",
        x"09",
        x"4C",
        x"B4",
        x"B5",
        x"B6",
        x"B5",
        x"BE",
        x"B4",
        x"B0",
        x"BF",
        x"C5",
        x"C2",
        x"B0",
        x"B0",
        x"83",
        x"81",
        x"0E",
        x"0A",
        x"CD",
        x"B4",
        x"B5",
        x"C3",
        x"C4",
        x"C2",
        x"BF",
        x"C9",
        x"B0",
        x"B5",
        x"BE",
        x"B5",
        x"BD",
        x"C9",
        x"B0",
        x"C4",
        x"B1",
        x"BE",
        x"BB",
        x"C3",
        x"13",
        x"0B",
        x"2A",
        x"BD",
        x"B9",
        x"C3",
        x"C3",
        x"B9",
        x"BF",
        x"BE",
        x"07",
        x"0A",
        x"67",
        x"FB",
        x"E0",
        x"F9",
        x"E4",
        x"E1",
        x"E5",
        x"F2",
        x"07",
        x"0A",
        x"67",
        x"EF",
        x"F7",
        x"F4",
        x"E0",
        x"F2",
        x"E5",
        x"F9",
        x"E1",
        x"EC",
        x"F0",
        x"0A",
        x"0A",
        x"89",
        x"E4",
        x"EE",
        x"F5",
        x"EF",
        x"F2",
        x"05",
        x"0A",
        x"11",
        x"C2",
        x"B5",
        x"B1",
        x"B4",
        x"C9",
        x"B0",
        x"CB",
        x"07",
        x"0A",
        x"58",
        x"C0",
        x"BC",
        x"B1",
        x"C9",
        x"B5",
        x"C2",
        x"B0",
        x"BF",
        x"BE",
        x"B5",
        x"0A",
        x"0A",
        x"96",
        x"C2",
        x"BF",
        x"C5",
        x"BE",
        x"B4",
        x"05",
        x"0A",
        x"6E",
        x"C4",
        x"C7",
        x"BF",
        x"03",
        x"09",
        x"B6",
        x"AC",
        x"B0",
        x"AD",
        x"AE",
        x"AF",
        x"DC",
        x"DD",
        x"DE",
        x"DF",
        x"B0",
        x"0C",
        x"0D",
        x"0E",
        x"0F",
        x"0E",
        x"0A",
        x"D6",
        x"B2",
        x"BF",
        x"BE",
        x"C5",
        x"C3",
        x"B0",
        x"C4",
        x"B1",
        x"BE",
        x"BB",
        x"B0",
        x"B6",
        x"BF",
        x"C2",
        x"B0",
        x"B0",
        x"A0",
        x"A0",
        x"A0",
        x"A0",
        x"B0",
        x"C0",
        x"C4",
        x"C3",
        x"18",
        x"0B",
        x"72",
        x"C0",
        x"C5",
        x"C3",
        x"B8",
        x"B0",
        x"C3",
        x"C4",
        x"B1",
        x"C2",
        x"C4",
        x"B0",
        x"B2",
        x"C5",
        x"C4",
        x"C4",
        x"BF",
        x"BE",
        x"11",
        x"0A",
        x"F0",
        x"B3",
        x"C2",
        x"B5",
        x"B4",
        x"B9",
        x"C4",
        x"06",
        x"0B",
        x"7F",
        x"B6",
        x"C2",
        x"B5",
        x"B5",
        x"B0",
        x"C0",
        x"BC",
        x"B1",
        x"C9",
        x"09",
        x"0B",
        x"7F",
        x"F0",
        x"F5",
        x"D2",
        x"E0",
        x"E0",
        x"E0",
        x"E5",
        x"F2",
        x"EF",
        x"E3",
        x"F3",
        x"E0",
        x"E8",
        x"E7",
        x"E9",
        x"E8",
        x"E0",
        x"E0",
        x"E0",
        x"F0",
        x"F5",
        x"D1",
        x"16",
        x"0B",
        x"5F",
        x"A1",
        x"C5",
        x"C0",
        x"B0",
        x"B0",
        x"B0",
        x"B8",
        x"B9",
        x"B7",
        x"B8",
        x"B0",
        x"C3",
        x"B3",
        x"BF",
        x"C2",
        x"B5",
        x"B0",
        x"B0",
        x"B0",
        x"A2",
        x"C5",
        x"C0",
        x"16",
        x"0B",
        x"40",
        x"F0",
        x"F5",
        x"D2",
        x"03",
        x"0B",
        x"5F",
        x"A2",
        x"C5",
        x"C0",
        x"03",
        x"08",
        x"E0",
        x"A1",
        x"C5",
        x"C0",
        x"03",
        x"0B",
        x"40",
        x"B0",
        x"B0",
        x"B0",
        x"03",
        x"0B",
        x"5F",
        x"B0",
        x"B0",
        x"B0",
        x"03",
        x"08",
        x"E0",
        x"B0",
        x"B0",
        x"B0",
        x"03",
        x"0B",
        x"40",
        x"AC",
        x"B0",
        x"BE",
        x"B1",
        x"BD",
        x"B3",
        x"BF",
        x"B0",
        x"BC",
        x"B9",
        x"BD",
        x"B9",
        x"C4",
        x"B5",
        x"B4",
        x"B0",
        x"A1",
        x"A9",
        x"A8",
        x"A0",
        x"14",
        x"0B",
        x"3B",
        x"C4",
        x"B1",
        x"BE",
        x"BB",
        x"04",
        x"0A",
        x"EC",
        x"BE",
        x"BF",
        x"C4",
        x"B8",
        x"B9",
        x"BE",
        x"B7",
        x"07",
        x"09",
        x"CA",
        x"A0",
        x"A0",
        x"A0",
        x"B0",
        x"B0",
        x"05",
        x"09",
        x"8A",
        x"B2",
        x"BF",
        x"BE",
        x"C5",
        x"C3",
        x"05",
        x"0A",
        x"EA",
        x"B6",
        x"C2",
        x"B5",
        x"B5",
        x"B0",
        x"C0",
        x"BC",
        x"B1",
        x"C9",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"B0",
        x"12",
        x"0A",
        x"E8",
        x"A2",
        x"B0",
        x"B3",
        x"C2",
        x"B5",
        x"B4",
        x"B9",
        x"C4",
        x"C3",
        x"09",
        x"09",
        x"C8",
        x"A1",
        x"B0",
        x"B3",
        x"C2",
        x"B5",
        x"B4",
        x"B9",
        x"C4",
        x"B0",
        x"09",
        x"09",
        x"C8",
        x"A2",
        x"B0",
        x"B3",
        x"BF",
        x"B9",
        x"BE",
        x"C3",
        x"B0",
        x"B0",
        x"09",
        x"0A",
        x"E8",
        x"A1",
        x"B0",
        x"B3",
        x"BF",
        x"B9",
        x"BE",
        x"B0",
        x"B0",
        x"B0",
        x"09",
        x"0A",
        x"E8",
        x"C5",
        x"C0",
        x"C2",
        x"B9",
        x"B7",
        x"B8",
        x"C4",
        x"07",
        x"0A",
        x"E6",
        x"C4",
        x"B1",
        x"B2",
        x"BC",
        x"B5",
        x"B0",
        x"B0",
        x"07",
        x"0A",
        x"E6"

    );
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";

begin
    process(clk)
    begin
        if rising_edge(clk) then
            if (oe_n = '0' and ce_n = '0') then
                data <= ROM(conv_integer(addr));
            end if;
        end if;
    end process;

end behavioral;