library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity IC7052 is
    port(
        clk  : in  std_logic;
        oe_n   : in  std_logic;
        ce_n   : in  std_logic;
        addr : in  std_logic_vector(7 downto 0);
        data : out std_logic_vector(3 downto 0)
    );
end IC7052;


--=INDEX($B$1:$B$256,ROWS(B1:$B$256))

architecture behavioral of IC7052 is
    type rom_type is array (255 downto 0) of std_logic_vector(3 downto 0);
    signal ROM : rom_type := (
        x"C",
        x"E",
        x"C",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"3",
        x"E",
        x"3",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"C",
        x"E",
        x"C",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"3",
        x"E",
        x"3",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"A",
        x"E",
        x"A",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"B",
        x"E",
        x"B",
        x"0",
        x"B",
        x"E",
        x"B",
        x"0",
        x"A",
        x"E",
        x"A",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"E",
        x"E",
        x"E",
        x"0",
        x"C",
        x"E",
        x"C",
        x"0",
        x"C",
        x"E",
        x"C",
        x"0",
        x"C",
        x"E",
        x"C",
        x"0",
        x"C",
        x"E",
        x"C",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"F",
        x"E",
        x"F",
        x"0",
        x"F",
        x"E",
        x"F",
        x"0",
        x"F",
        x"E",
        x"F",
        x"0",
        x"F",
        x"E",
        x"F",
        x"0",
        x"3",
        x"E",
        x"3",
        x"0",
        x"3",
        x"E",
        x"3",
        x"0",
        x"3",
        x"E",
        x"3",
        x"0",
        x"3",
        x"E",
        x"3",
        x"0",
        x"F",
        x"E",
        x"F",
        x"0",
        x"7",
        x"E",
        x"7",
        x"0",
        x"3",
        x"E",
        x"3",
        x"0",
        x"5",
        x"0",
        x"5",
        x"0",
        x"3",
        x"E",
        x"3",
        x"0",
        x"2",
        x"E",
        x"2",
        x"0",
        x"2",
        x"E",
        x"2",
        x"0",
        x"2",
        x"E",
        x"2",
        x"0");
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";

begin
    process(clk)
    begin
        if rising_edge(clk) then
            if (oe_n = '0' and ce_n = '0') then
                data <= ROM(conv_integer(addr));
            end if;
        end if;
    end process;

end behavioral;