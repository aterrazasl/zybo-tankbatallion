library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity M2716 is
    port(
        clk  : in  std_logic;
        oe_n   : in  std_logic;
        ce_n   : in  std_logic;
        addr : in  std_logic_vector(10 downto 0);
        data : out std_logic_vector(7 downto 0)
    );
end M2716;

architecture behavioral of M2716 is
    type rom_type is array (2047 downto 0) of std_logic_vector(7 downto 0);
    signal ROM : rom_type := (
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"F8",
        x"F8",
        x"52",
        x"5E",
        x"52",
        x"F8",
        x"F8",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"06",
        x"0F",
        x"59",
        x"51",
        x"03",
        x"02",
        x"00",
        x"00",
        x"00",
        x"00",
        x"07",
        x"5F",
        x"5F",
        x"00",
        x"00",
        x"00",
        x"43",
        x"47",
        x"4F",
        x"5D",
        x"79",
        x"71",
        x"61",
        x"00",
        x"07",
        x"0F",
        x"78",
        x"78",
        x"0F",
        x"07",
        x"00",
        x"00",
        x"63",
        x"77",
        x"3E",
        x"1C",
        x"3E",
        x"77",
        x"63",
        x"00",
        x"7F",
        x"7F",
        x"38",
        x"1C",
        x"38",
        x"7F",
        x"7F",
        x"00",
        x"0F",
        x"1F",
        x"38",
        x"70",
        x"38",
        x"1F",
        x"0F",
        x"00",
        x"3F",
        x"7F",
        x"40",
        x"40",
        x"40",
        x"7F",
        x"3F",
        x"00",
        x"01",
        x"01",
        x"7F",
        x"7F",
        x"01",
        x"01",
        x"00",
        x"00",
        x"30",
        x"7A",
        x"4B",
        x"49",
        x"49",
        x"6F",
        x"26",
        x"00",
        x"4E",
        x"6F",
        x"79",
        x"31",
        x"11",
        x"7F",
        x"7F",
        x"00",
        x"5E",
        x"3F",
        x"71",
        x"51",
        x"41",
        x"7F",
        x"3E",
        x"00",
        x"0E",
        x"1F",
        x"11",
        x"11",
        x"11",
        x"7F",
        x"7F",
        x"00",
        x"3E",
        x"7F",
        x"41",
        x"41",
        x"41",
        x"7F",
        x"3E",
        x"00",
        x"7F",
        x"7F",
        x"38",
        x"1C",
        x"0E",
        x"7F",
        x"7F",
        x"00",
        x"7F",
        x"7F",
        x"0E",
        x"1C",
        x"0E",
        x"7F",
        x"7F",
        x"00",
        x"40",
        x"40",
        x"40",
        x"40",
        x"7F",
        x"7F",
        x"00",
        x"00",
        x"FF",
        x"01",
        x"01",
        x"01",
        x"01",
        x"01",
        x"01",
        x"01",
        x"FF",
        x"80",
        x"80",
        x"80",
        x"80",
        x"80",
        x"80",
        x"80",
        x"41",
        x"41",
        x"7F",
        x"7F",
        x"41",
        x"41",
        x"00",
        x"00",
        x"7F",
        x"7F",
        x"08",
        x"08",
        x"08",
        x"7F",
        x"7F",
        x"00",
        x"79",
        x"79",
        x"49",
        x"41",
        x"63",
        x"3E",
        x"1C",
        x"00",
        x"01",
        x"09",
        x"09",
        x"09",
        x"09",
        x"7F",
        x"7F",
        x"00",
        x"41",
        x"49",
        x"49",
        x"49",
        x"7F",
        x"7F",
        x"00",
        x"00",
        x"1C",
        x"3E",
        x"63",
        x"41",
        x"41",
        x"7F",
        x"7F",
        x"00",
        x"22",
        x"63",
        x"41",
        x"41",
        x"63",
        x"3E",
        x"1C",
        x"00",
        x"36",
        x"7F",
        x"49",
        x"49",
        x"49",
        x"7F",
        x"7F",
        x"00",
        x"7C",
        x"7E",
        x"13",
        x"11",
        x"13",
        x"7E",
        x"7C",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"C3",
        x"C3",
        x"C3",
        x"C3",
        x"FF",
        x"7E",
        x"00",
        x"00",
        x"C3",
        x"C3",
        x"C3",
        x"00",
        x"00",
        x"7E",
        x"FF",
        x"C3",
        x"7F",
        x"00",
        x"00",
        x"7E",
        x"FF",
        x"C3",
        x"C3",
        x"C3",
        x"FF",
        x"C0",
        x"C0",
        x"FF",
        x"FF",
        x"C0",
        x"C0",
        x"FF",
        x"01",
        x"01",
        x"01",
        x"01",
        x"01",
        x"01",
        x"01",
        x"FF",
        x"80",
        x"80",
        x"80",
        x"80",
        x"80",
        x"80",
        x"80",
        x"FF",
        x"1E",
        x"3F",
        x"69",
        x"49",
        x"49",
        x"4F",
        x"06",
        x"00",
        x"30",
        x"76",
        x"59",
        x"59",
        x"4D",
        x"4F",
        x"36",
        x"00",
        x"03",
        x"07",
        x"0D",
        x"79",
        x"71",
        x"03",
        x"03",
        x"00",
        x"30",
        x"79",
        x"49",
        x"49",
        x"4B",
        x"7E",
        x"3C",
        x"00",
        x"38",
        x"7D",
        x"45",
        x"45",
        x"45",
        x"67",
        x"27",
        x"00",
        x"10",
        x"7F",
        x"7F",
        x"13",
        x"16",
        x"1C",
        x"18",
        x"00",
        x"31",
        x"7B",
        x"4F",
        x"4D",
        x"49",
        x"61",
        x"20",
        x"00",
        x"46",
        x"4F",
        x"5D",
        x"59",
        x"79",
        x"73",
        x"62",
        x"00",
        x"40",
        x"40",
        x"7F",
        x"7F",
        x"42",
        x"40",
        x"00",
        x"00",
        x"1C",
        x"3E",
        x"43",
        x"41",
        x"61",
        x"3E",
        x"1C",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"1F",
        x"1F",
        x"4A",
        x"7A",
        x"4A",
        x"1F",
        x"1F",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"40",
        x"C0",
        x"8A",
        x"9A",
        x"F0",
        x"60",
        x"00",
        x"00",
        x"00",
        x"FA",
        x"FA",
        x"E0",
        x"00",
        x"00",
        x"00",
        x"86",
        x"8E",
        x"9E",
        x"BA",
        x"F2",
        x"E2",
        x"C2",
        x"00",
        x"00",
        x"E0",
        x"F0",
        x"1E",
        x"1E",
        x"F0",
        x"E0",
        x"00",
        x"C6",
        x"EE",
        x"7C",
        x"38",
        x"7C",
        x"EE",
        x"C6",
        x"00",
        x"FE",
        x"FE",
        x"1C",
        x"38",
        x"1C",
        x"FE",
        x"FE",
        x"00",
        x"F0",
        x"F8",
        x"1C",
        x"0E",
        x"1C",
        x"F8",
        x"F0",
        x"00",
        x"FC",
        x"FE",
        x"02",
        x"02",
        x"02",
        x"FE",
        x"FC",
        x"00",
        x"00",
        x"80",
        x"80",
        x"FE",
        x"FE",
        x"80",
        x"80",
        x"00",
        x"64",
        x"F6",
        x"92",
        x"92",
        x"D2",
        x"5E",
        x"0C",
        x"00",
        x"FE",
        x"FE",
        x"88",
        x"8C",
        x"9E",
        x"F6",
        x"72",
        x"00",
        x"7C",
        x"FE",
        x"82",
        x"8A",
        x"8E",
        x"FC",
        x"7A",
        x"00",
        x"FE",
        x"FE",
        x"88",
        x"88",
        x"88",
        x"F8",
        x"70",
        x"00",
        x"7C",
        x"FE",
        x"82",
        x"82",
        x"82",
        x"FE",
        x"7C",
        x"00",
        x"FE",
        x"FE",
        x"70",
        x"38",
        x"1C",
        x"FE",
        x"FE",
        x"00",
        x"FE",
        x"FE",
        x"70",
        x"38",
        x"70",
        x"FE",
        x"FE",
        x"00",
        x"00",
        x"FE",
        x"FE",
        x"02",
        x"02",
        x"02",
        x"02",
        x"00",
        x"FE",
        x"FE",
        x"18",
        x"3C",
        x"6E",
        x"C6",
        x"82",
        x"00",
        x"04",
        x"06",
        x"02",
        x"02",
        x"02",
        x"FE",
        x"FC",
        x"00",
        x"00",
        x"82",
        x"82",
        x"FE",
        x"FE",
        x"82",
        x"82",
        x"00",
        x"FE",
        x"FE",
        x"10",
        x"10",
        x"10",
        x"FE",
        x"FE",
        x"00",
        x"38",
        x"7C",
        x"C6",
        x"82",
        x"92",
        x"9E",
        x"9E",
        x"00",
        x"FE",
        x"FE",
        x"90",
        x"90",
        x"90",
        x"90",
        x"80",
        x"00",
        x"00",
        x"FE",
        x"FE",
        x"92",
        x"92",
        x"92",
        x"82",
        x"00",
        x"FE",
        x"FE",
        x"82",
        x"82",
        x"C6",
        x"7C",
        x"38",
        x"00",
        x"38",
        x"7C",
        x"C6",
        x"82",
        x"82",
        x"C6",
        x"44",
        x"00",
        x"FE",
        x"FE",
        x"92",
        x"92",
        x"92",
        x"FE",
        x"6C",
        x"00",
        x"3E",
        x"7E",
        x"C8",
        x"88",
        x"C8",
        x"7E",
        x"3E",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"DB",
        x"DB",
        x"FF",
        x"FF",
        x"7F",
        x"00",
        x"00",
        x"FF",
        x"FF",
        x"7F",
        x"00",
        x"00",
        x"1F",
        x"DF",
        x"DB",
        x"DB",
        x"00",
        x"00",
        x"FF",
        x"FF",
        x"C0",
        x"C0",
        x"C0",
        x"C0",
        x"3C",
        x"42",
        x"99",
        x"A5",
        x"A5",
        x"81",
        x"42",
        x"3C",
        x"00",
        x"FE",
        x"FE",
        x"92",
        x"92",
        x"92",
        x"FE",
        x"6C",
        x"00",
        x"60",
        x"E0",
        x"CA",
        x"CA",
        x"DA",
        x"F0",
        x"60",
        x"00",
        x"60",
        x"F2",
        x"92",
        x"92",
        x"96",
        x"FC",
        x"78",
        x"00",
        x"6C",
        x"F2",
        x"B2",
        x"9A",
        x"9A",
        x"6E",
        x"0C",
        x"00",
        x"C0",
        x"C0",
        x"8E",
        x"9E",
        x"B0",
        x"E0",
        x"C0",
        x"00",
        x"3C",
        x"7E",
        x"D2",
        x"92",
        x"92",
        x"9E",
        x"0C",
        x"00",
        x"E4",
        x"E6",
        x"A2",
        x"A2",
        x"A2",
        x"BE",
        x"1C",
        x"00",
        x"18",
        x"38",
        x"68",
        x"C8",
        x"FE",
        x"FE",
        x"08",
        x"00",
        x"04",
        x"86",
        x"92",
        x"B2",
        x"F2",
        x"DE",
        x"8C",
        x"00",
        x"46",
        x"CE",
        x"9E",
        x"9A",
        x"BA",
        x"F2",
        x"62",
        x"00",
        x"00",
        x"02",
        x"42",
        x"FE",
        x"FE",
        x"02",
        x"02",
        x"00",
        x"38",
        x"7C",
        x"86",
        x"82",
        x"C2",
        x"7C",
        x"38",
        x"80",
        x"C0",
        x"E0",
        x"E0",
        x"F0",
        x"F0",
        x"F8",
        x"F8",
        x"00",
        x"00",
        x"01",
        x"01",
        x"03",
        x"03",
        x"07",
        x"07",
        x"8C",
        x"84",
        x"34",
        x"74",
        x"76",
        x"06",
        x"06",
        x"FE",
        x"0C",
        x"0C",
        x"0C",
        x"0E",
        x"1F",
        x"1C",
        x"1C",
        x"1F",
        x"FE",
        x"FE",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"FF",
        x"FF",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"2A",
        x"BE",
        x"FC",
        x"B8",
        x"60",
        x"E0",
        x"C8",
        x"F4",
        x"00",
        x"00",
        x"03",
        x"07",
        x"67",
        x"67",
        x"32",
        x"7F",
        x"FC",
        x"C4",
        x"E0",
        x"60",
        x"B8",
        x"FC",
        x"BE",
        x"2A",
        x"7F",
        x"32",
        x"67",
        x"67",
        x"07",
        x"03",
        x"00",
        x"00",
        x"F8",
        x"38",
        x"38",
        x"F8",
        x"70",
        x"30",
        x"30",
        x"B0",
        x"7F",
        x"60",
        x"60",
        x"6E",
        x"2E",
        x"2C",
        x"21",
        x"31",
        x"E0",
        x"E0",
        x"C0",
        x"C0",
        x"80",
        x"80",
        x"00",
        x"00",
        x"1F",
        x"1F",
        x"0F",
        x"0F",
        x"07",
        x"07",
        x"03",
        x"01",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"FF",
        x"FF",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"7F",
        x"7F",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"C0",
        x"E0",
        x"E6",
        x"E6",
        x"4C",
        x"FE",
        x"54",
        x"7D",
        x"3F",
        x"1D",
        x"06",
        x"07",
        x"23",
        x"3F",
        x"FE",
        x"4C",
        x"E6",
        x"E6",
        x"E0",
        x"C0",
        x"00",
        x"00",
        x"2F",
        x"13",
        x"07",
        x"06",
        x"1D",
        x"3F",
        x"7D",
        x"54",
        x"00",
        x"00",
        x"80",
        x"C0",
        x"C0",
        x"C0",
        x"E0",
        x"F0",
        x"00",
        x"06",
        x"1F",
        x"01",
        x"07",
        x"03",
        x"03",
        x"07",
        x"F8",
        x"F0",
        x"EC",
        x"98",
        x"60",
        x"C0",
        x"00",
        x"00",
        x"1F",
        x"0F",
        x"0F",
        x"07",
        x"04",
        x"01",
        x"FF",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"39",
        x"49",
        x"49",
        x"3E",
        x"00",
        x"7F",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"36",
        x"49",
        x"49",
        x"49",
        x"36",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"31",
        x"4B",
        x"45",
        x"41",
        x"21",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"39",
        x"45",
        x"45",
        x"45",
        x"27",
        x"00",
        x"40",
        x"7F",
        x"42",
        x"00",
        x"00",
        x"00",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"30",
        x"49",
        x"49",
        x"4A",
        x"3C",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"3E",
        x"41",
        x"41",
        x"41",
        x"3E",
        x"00",
        x"31",
        x"4B",
        x"45",
        x"41",
        x"21",
        x"00",
        x"00",
        x"00",
        x"FF",
        x"80",
        x"20",
        x"E0",
        x"F0",
        x"F0",
        x"F8",
        x"00",
        x"00",
        x"03",
        x"06",
        x"19",
        x"37",
        x"0F",
        x"1F",
        x"E0",
        x"C0",
        x"C0",
        x"E0",
        x"80",
        x"F8",
        x"60",
        x"00",
        x"0F",
        x"07",
        x"03",
        x"03",
        x"03",
        x"01",
        x"00",
        x"00",
        x"FE",
        x"00",
        x"7C",
        x"92",
        x"92",
        x"9C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"7C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"7C",
        x"6C",
        x"92",
        x"92",
        x"92",
        x"6C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"7C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"7C",
        x"00",
        x"84",
        x"82",
        x"A2",
        x"D2",
        x"8C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"7C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"7C",
        x"00",
        x"00",
        x"42",
        x"FE",
        x"02",
        x"00",
        x"E4",
        x"A2",
        x"A2",
        x"A2",
        x"9C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"7C",
        x"00",
        x"00",
        x"00",
        x"3C",
        x"52",
        x"92",
        x"92",
        x"0C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"82",
        x"7C",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"84",
        x"82",
        x"A2",
        x"D2",
        x"8C",
        x"00",
        x"7C",
        x"82",
        x"82",
        x"82",
        x"7C",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"FC",
        x"FC",
        x"FC",
        x"C0",
        x"60",
        x"30",
        x"00",
        x"00",
        x"0F",
        x"0F",
        x"0F",
        x"03",
        x"06",
        x"64",
        x"18",
        x"30",
        x"60",
        x"C0",
        x"FC",
        x"FC",
        x"FC",
        x"00",
        x"7C",
        x"64",
        x"06",
        x"03",
        x"0F",
        x"0F",
        x"0F",
        x"00",
        x"00",
        x"00",
        x"E0",
        x"E0",
        x"E0",
        x"80",
        x"C0",
        x"4C",
        x"00",
        x"00",
        x"7F",
        x"7F",
        x"7F",
        x"07",
        x"0C",
        x"18",
        x"7C",
        x"4C",
        x"C0",
        x"80",
        x"E0",
        x"E0",
        x"E0",
        x"00",
        x"30",
        x"18",
        x"0C",
        x"07",
        x"7F",
        x"7F",
        x"7F",
        x"00",
        x"00",
        x"00",
        x"80",
        x"80",
        x"00",
        x"1C",
        x"DC",
        x"7C",
        x"00",
        x"00",
        x"03",
        x"03",
        x"01",
        x"71",
        x"77",
        x"7C",
        x"3C",
        x"3C",
        x"7C",
        x"DC",
        x"9C",
        x"1C",
        x"1C",
        x"00",
        x"78",
        x"78",
        x"7C",
        x"76",
        x"73",
        x"71",
        x"70",
        x"00",
        x"00",
        x"00",
        x"1C",
        x"1C",
        x"9C",
        x"DC",
        x"7C",
        x"3C",
        x"00",
        x"00",
        x"70",
        x"71",
        x"73",
        x"76",
        x"7C",
        x"78",
        x"3C",
        x"7C",
        x"DC",
        x"1C",
        x"00",
        x"80",
        x"80",
        x"00",
        x"78",
        x"7C",
        x"77",
        x"71",
        x"01",
        x"03",
        x"03",
        x"00",
        x"00",
        x"00",
        x"FC",
        x"FC",
        x"FC",
        x"F0",
        x"F8",
        x"F8",
        x"00",
        x"00",
        x"03",
        x"03",
        x"03",
        x"00",
        x"01",
        x"63",
        x"F8",
        x"F8",
        x"F8",
        x"F0",
        x"FC",
        x"FC",
        x"FC",
        x"00",
        x"7F",
        x"63",
        x"01",
        x"00",
        x"03",
        x"03",
        x"03",
        x"00",
        x"00",
        x"00",
        x"80",
        x"80",
        x"80",
        x"00",
        x"00",
        x"8C",
        x"00",
        x"00",
        x"7F",
        x"7F",
        x"7F",
        x"1E",
        x"3F",
        x"3F",
        x"FC",
        x"8C",
        x"00",
        x"00",
        x"80",
        x"80",
        x"80",
        x"00",
        x"3F",
        x"3F",
        x"3F",
        x"1E",
        x"7F",
        x"7F",
        x"7F",
        x"00",
        x"00",
        x"00",
        x"80",
        x"80",
        x"00",
        x"00",
        x"00",
        x"9C",
        x"00",
        x"00",
        x"03",
        x"03",
        x"01",
        x"01",
        x"01",
        x"73",
        x"DC",
        x"FC",
        x"FC",
        x"FC",
        x"FC",
        x"DC",
        x"1C",
        x"00",
        x"77",
        x"7F",
        x"7F",
        x"7F",
        x"7F",
        x"77",
        x"70",
        x"00",
        x"00",
        x"00",
        x"1C",
        x"DC",
        x"FC",
        x"FC",
        x"FC",
        x"FC",
        x"00",
        x"00",
        x"70",
        x"77",
        x"7F",
        x"7F",
        x"7F",
        x"7F",
        x"DC",
        x"9C",
        x"00",
        x"00",
        x"00",
        x"80",
        x"80",
        x"00",
        x"77",
        x"73",
        x"01",
        x"01",
        x"01",
        x"03",
        x"03",
        x"00",
        x"80",
        x"48",
        x"28",
        x"13",
        x"27",
        x"0F",
        x"0F",
        x"0E",
        x"50",
        x"48",
        x"3D",
        x"83",
        x"9F",
        x"DE",
        x"FF",
        x"3F",
        x"74",
        x"FF",
        x"CB",
        x"B5",
        x"7F",
        x"FF",
        x"FE",
        x"CF",
        x"01",
        x"0A",
        x"94",
        x"84",
        x"F0",
        x"3C",
        x"DE",
        x"EF",
        x"0D",
        x"07",
        x"6F",
        x"FF",
        x"FB",
        x"FF",
        x"EF",
        x"7F",
        x"BF",
        x"FF",
        x"FD",
        x"9C",
        x"C1",
        x"61",
        x"AD",
        x"E7",
        x"B7",
        x"FF",
        x"FB",
        x"67",
        x"0F",
        x"2F",
        x"D8",
        x"87",
        x"F7",
        x"FB",
        x"F7",
        x"FA",
        x"F7",
        x"EF",
        x"7F",
        x"FF",
        x"5D",
        x"1B",
        x"1B",
        x"3D",
        x"3F",
        x"19",
        x"06",
        x"0F",
        x"83",
        x"E1",
        x"ED",
        x"D3",
        x"C5",
        x"DC",
        x"7D",
        x"BF",
        x"EF",
        x"8B",
        x"5D",
        x"2F",
        x"17",
        x"CB",
        x"EF",
        x"FF",
        x"FF",
        x"F8",
        x"DE",
        x"EF",
        x"F7",
        x"F6",
        x"EE",
        x"FE",
        x"0F",
        x"03",
        x"13",
        x"19",
        x"30",
        x"62",
        x"C4",
        x"80",
        x"FF",
        x"FF",
        x"DF",
        x"F7",
        x"DE",
        x"0F",
        x"00",
        x"00",
        x"FF",
        x"FF",
        x"FE",
        x"6D",
        x"73",
        x"7F",
        x"1E",
        x"00",
        x"FC",
        x"58",
        x"C0",
        x"C8",
        x"98",
        x"0C",
        x"02",
        x"00",
        x"00",
        x"20",
        x"20",
        x"10",
        x"09",
        x"0D",
        x"02",
        x"04",
        x"00",
        x"20",
        x"20",
        x"4E",
        x"1F",
        x"39",
        x"36",
        x"6F",
        x"00",
        x"00",
        x"04",
        x"E2",
        x"F8",
        x"7C",
        x"BC",
        x"FA",
        x"00",
        x"00",
        x"04",
        x"48",
        x"90",
        x"A0",
        x"40",
        x"30",
        x"00",
        x"03",
        x"0F",
        x"1D",
        x"1E",
        x"0D",
        x"1B",
        x"1D",
        x"FF",
        x"6D",
        x"B6",
        x"FE",
        x"E6",
        x"E8",
        x"F6",
        x"7B",
        x"E7",
        x"FF",
        x"DF",
        x"F3",
        x"A7",
        x"17",
        x"AF",
        x"CF",
        x"80",
        x"C0",
        x"61",
        x"B6",
        x"B4",
        x"66",
        x"F4",
        x"B0",
        x"1B",
        x"0F",
        x"07",
        x"01",
        x"11",
        x"09",
        x"04",
        x"04",
        x"D7",
        x"F1",
        x"6D",
        x"FD",
        x"FE",
        x"FE",
        x"DB",
        x"67",
        x"E3",
        x"4F",
        x"2F",
        x"77",
        x"7F",
        x"FE",
        x"FD",
        x"AB",
        x"C0",
        x"E0",
        x"60",
        x"B0",
        x"F0",
        x"E4",
        x"08",
        x"00",
        x"03",
        x"0D",
        x"09",
        x"18",
        x"30",
        x"20",
        x"00",
        x"00",
        x"7F",
        x"1C",
        x"00",
        x"24",
        x"38",
        x"28",
        x"00",
        x"00",
        x"D6",
        x"FE",
        x"78",
        x"02",
        x"08",
        x"00",
        x"00",
        x"00",
        x"C0",
        x"A0",
        x"10",
        x"08",
        x"04",
        x"04",
        x"00",
        x"00",
        x"B3",
        x"B6",
        x"DC",
        x"F9",
        x"F0",
        x"5E",
        x"3C",
        x"B8",
        x"9C",
        x"C0",
        x"64",
        x"7F",
        x"BB",
        x"DF",
        x"19",
        x"FC",
        x"BF",
        x"10",
        x"69",
        x"FD",
        x"DD",
        x"8C",
        x"86",
        x"53",
        x"75",
        x"38",
        x"9D",
        x"97",
        x"3F",
        x"79",
        x"64",
        x"8E",
        x"00",
        x"02",
        x"66",
        x"6C",
        x"F8",
        x"EC",
        x"38",
        x"78",
        x"00",
        x"60",
        x"32",
        x"1F",
        x"0B",
        x"1D",
        x"1F",
        x"0E",
        x"30",
        x"38",
        x"7C",
        x"C8",
        x"FC",
        x"4E",
        x"02",
        x"00",
        x"7C",
        x"0E",
        x"0B",
        x"1D",
        x"1F",
        x"3B",
        x"70",
        x"40",
        x"00",
        x"00",
        x"00",
        x"44",
        x"E8",
        x"B8",
        x"F0",
        x"60",
        x"00",
        x"00",
        x"00",
        x"04",
        x"32",
        x"1F",
        x"0D",
        x"06",
        x"30",
        x"78",
        x"E0",
        x"70",
        x"50",
        x"08",
        x"00",
        x"00",
        x"1E",
        x"09",
        x"1F",
        x"3B",
        x"22",
        x"02",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"55",
        x"AA",
        x"55",
        x"AA",
        x"55",
        x"AA",
        x"55",
        x"AA",
        x"00",
        x"38",
        x"7C",
        x"86",
        x"82",
        x"C2",
        x"7C",
        x"38",
        x"00",
        x"6C",
        x"F2",
        x"B2",
        x"9A",
        x"9A",
        x"6E",
        x"0C",
        x"00",
        x"60",
        x"F2",
        x"92",
        x"92",
        x"96",
        x"FC",
        x"78",
        x"00",
        x"00",
        x"02",
        x"42",
        x"FE",
        x"FE",
        x"02",
        x"02",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"0E",
        x"0E",
        x"0E",
        x"0E",
        x"00",
        x"00",
        x"00",
        x"00",
        x"E0",
        x"E0",
        x"00",
        x"E0",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"0E",
        x"0E",
        x"00",
        x"0E",
        x"00",
        x"00",
        x"00",
        x"00",
        x"E0",
        x"E0",
        x"E0",
        x"E0",
        x"E0",
        x"E0",
        x"00",
        x"E0",
        x"E0",
        x"E0",
        x"E0",
        x"E0",
        x"0E",
        x"0E",
        x"0E",
        x"0E",
        x"0E",
        x"0E",
        x"00",
        x"0E",
        x"EE",
        x"EE",
        x"0E",
        x"EE",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"EE",
        x"EE",
        x"E0",
        x"EE",
        x"EE",
        x"EE",
        x"0E",
        x"EE",
        x"EE",
        x"EE",
        x"E0",
        x"EE",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00",
        x"00");
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";

begin
    process(clk)
    begin
        if rising_edge(clk) then
            if (oe_n = '0' and ce_n = '0') then
                data <= ROM(conv_integer(addr));
            end if;
        end if;
    end process;

end behavioral;